��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�Xx�(c���J3v����=�I��O&��2��O�j
m�ҡ��rz�z�v	R��"�R��췰Z�ʁ�����,�>�����P��$�Y��B}�R�w�Y�["3̊���e�Hʩ�D�$���s2�l*���)f�|}3���K�q s�])a�'�<7�������0ꐿ�	�O���K�"BH8>�?�ψ��ޥ���Hd�I-�m3v	G�W=U5}��JMi=���KR5��꯼p	7���{����z��) ����lʉgv���:rf�m{v��9�3�B"���Ԩ����+�p-2�9ᔚ��Ao�J�T{���i8p]E�sd:�R�����Iv��t��s���}�'��bR2m,� �Kɾ帢���N%3gv�cٮy&��"\��m�ia�J���|_�������y�����]&L�]Ш["��|�
���Pk`�e�,'8M�X��|��4��g�	;N��P�D���i6�M:Ǔ�\
Է�l7�4ݫ�ZEܧ���k+;>��j�K"���1�6�G�^Z���.a������7/��C�v�~��yz�e4:�e�v����6� ������6��B�,��`[�"	"J�E�L��SYC�|rͽ��Jqa���3��5CO�M�i�f1x��g?�O�OR��xFF�⤻�j��B�f�
�kJ���&-)O�,�g���+K�h��1S��P�=2Q���w�����y,����a��&�A"~��k��<dmg�*/��1B�>c���g!4?��d,���9.m���_�H��lz�N�6N��~�	��K�6o�`����'<���9��$V��,|�0b+���t����b�!:BNGc�-{������	.����F��N>�ʐYN#�� ��
�y�%�YQ�V�d ��V��>c�G�v��<��4ۭ�n�~��,�gxK���U'�"خ��s�(�p}��{�8/N���@�X�BԨ:i�$zy�$���2����d+;��]h��P� gz�q|b�����!`^%�ΪIw����bK�2�,�ٙ���/�?w���eՀ�m1����ʧc�g�V*.��хF�B��;�$`�C�I��n�-ۓW4(U��Y�`��"�cɗ���0A;�6�H O�O��]/[3,
�(�H}d��3Ngb�!/7=遜��U~�+ء�Y���y*�vp�I��H۪�\%�4W6�jM���ay����m�g�I��t `�8�ݚ��՗!�^�!�i�V�+�|�h��5on�q�U�(?�\� ��M���?$*�*����")T_��j��ŕV�`W�K�R�]�Z$�G�AR^��E�����39̛��Y�)�_&�mi+,�J�ZrG�HJň龒��}���f$^�,f� '����04[Q���m��`��Հ0Pd�ruc�'w:�a3ɇ��	�4�ZX�_?d���IJQwdu�nD����`r����E1�O�s���dT܅�SDe�҆,�{�����������W1�L�-k�b=t��`�i��9�MK�U(_� �ZE�#Z@�܂Dx�;'�(�V_�?��u�n�� H��9�8�x��Nep?^�TV��!4�η[���e�qz�Z�WD�L�%MQd������ȧ� E7zO0nH�}�A�C�p?�ܪ@0��AF����Gb��EZ�����x-���i߬�偐_99]+l�)d�-�o���e���ܹ�S��=;0��	�nvѩ�ti)����xYW���휺������PǗ7TYb̺I_��i3Q�"�2�i�<{�X5�V����@\[�#R��8��j+U��*�OE�� H�ߓw��N����J6Oa۽�KC��a$��N���CC�<�B�ʡ�\`L��RVW�/k�q��⷟��oV��؇�\��H�i�(_uW�M��f�!>�}�X7B��аܢ(S#�%��c�V1�T�a`����Í[\� x 6tL���VYͱ�1t�%��S0�����͔.>/a������T�����Y��ڲpnY�X����N��/��Łơh��4��k��Z�t�'�Ι����B����ܥ���RF�ɿ�Nڰ*����F�#tJrZ��裣���B�F*�w;�u�p��"��&�U��˫����
=O�H$)�NX'z���8s!����������YΡ^�<켜�焵��a��3��2>�(�|LH8�/��|���ؑ�Zʲj�c�r���������'��'j?'R:�U�����i�ކ�4銛CB������b�.wЩ�g=;��Ϲ��X�</q�"��W�$J����+����4�$�T+G9�1�Q��V��}_7G=��Uf9�M�V2噢�����,@(?>9��].=������P�U���Kx�U���<1W��)�?���mH��᫾$������ ,}X�.��rɀz=���$�N��>����^J3[NZ�7C�͐ǈT{�wE-�:>0�lxG�`��ϰ�����lQ#��B�L�&"i�K.)c����˦^)b��������r�TC�H���z<؞0�2$�1fO{,���/g-8�^��X�eS���ʈ��re��kx��j��P	����Ꮋ�咄#ln�D��p�:����:���x�/Hд��D.���L&���R5��y����I��WZV�³}@�"�t�e��o$O�NO���Q� \(�i��gk3�x��͌�/#��Ur��0���� �\����,ֵ��O�$",G?COK�%U5�^c{�}qS�2�Q�ΉR� S�5����pV/K'�Q��M/S���qTgS?[Tآ�z�G�t�̾X��{K�b�
���yw-G(�}�<���AE���:h�~[����Ӄ�B�9��l��S��1ܫ�`�J��j}ٔ���u����o��g;�]�K����_�h%J^��V E��GH��+�d��#gu�~rxSWU������8bI�������sH�*��1I�3U��k���8����?���^!#������W:�D�1��.�:�Tpr lz�������"�Tdj��.u�]�� �,[|e�و���ݎ�S�[y�������od�>,����t�=p�a��s���"�7�������=iX��:"���ϗ��p���mNN�tl�n��s�e����񞂮�*t��ҩ��3�P�dβ^ڹ�����?�~����?LJ�3^Q6�e&�����P���
2��TD��Ĭ�Sj�L���h�����L���n���h+㧨��
�k�3�E�D�np�MU��)����W�H-4�����GsI��~y_�������c ��5Қ\�a^@���q7����~�����-݇Z�GCm�i�Ӓ�+h���SfR�iEA�5���ʿM��Q"�:��c	�;�  ^¿�y��J�FNɁG���fČ
�Eb��,�%m-�h���� Xk������u��imZ�lb'\���-^�e3vk[���U�TW�+H�d��]T���_��5���N�j
�{<a�i�>(���!���������myچ0;:c���Q��
��^%r�`��t��5U���|��ΰ�_Ͱ� �YaG{�U�v�����o|�������u�%�j���:eZ��d�������2~ޅ{�o�H���P����'!汮O�/#9o��{�1n S��x����D='�2��+���-�Ku��ysƷ�B&�����Ǟ���B���e�e3��o�Z26�ylQ n?".蝠��z��;z�u4Q}�g|����g��O۠A%\�������R��9�գ��2{���|繄|���|�YqK����i�+2��aI	��w����H���U�������+�*oG�J�������(�6ɳ��)ՃH�FeR$��TUMKJ��`ťO��;����4�
+�׉K�~'kv�ґz��?�!�ı���{��Q��1:�۰���j���K��ܯe�\��Xx�栂�EQ����/�h~g.�t�Ax(�>�3��s�l��S������^}�q�grT;6�#e)�I�]b�9Q���P�Ԋ���/6s���C��^ۅ�w����T�>�ч},�]̲[�̀��`����7.�G�� @��?�{h��+˝�O:d~o�TVB��zT�[:R���&��Z�V�k�'�Ů�ŋTh���6fOw�;�L!��U��W��'��\��|\��_/u49����>�j����#m��)L���m��҅�4 �^�|>()ߐN� �W�l/^����f���%+p:�}��/����I�'Hpo��-U�ݽz9�f�?+�#�����}s�^��~LDb�ZB�=���(*#ժ��6�IO|�� Z����;@Kzd�DԂ��v���`���ϰ�$�+�_�n�����6).��8�Q����g\�Q�����]/�A�N4�ۆZ.�YH	��P7�y�f�i��%�G�tS�Fі����d_=Kߐ}v���b&2��RH�b�Ҵb�cӧ�(�,�;-�̊���t�g�ٚc��
���u���:D�]I����|oq���c*@M����;	���j��B���3�{���C*���0j/���KZ�Vy#��!&����L��o2W� {"	�"�JĊJ�'�@ߢ��]M5���c��G3��HFӜ���/�e	ܸ��ɻ\8Ңrl]��o��`Hx�7��I>U�@�U��K+�Ey4eڦ�k�������tr�iw8��_8� o��ZGPO��Z��1�׽V�J��ޔ>C/E2�ۄِi�;�����AP�����k��ʐ@�?a�~��$w�|:t���}
NXTR�7$K���wY�_y�/.� )�^i�b��9�C�X�����{
%�|4?���&���=,3q�2]���T����>-��ND�=Y=+�f_������2;�UqCN/q7�z���]�*ea�x�PZD��"���"+1�('J0�M�_���j��w��*#M1Zc�PR�{3S!��VJKz��U�/�,]Pl�UϜ.1EԆ�����ۡf]��>����>��B�?z�v�/����@�ڝC}����5d-U�UG�P��+���]�?�3� ?0oh�����SH��]�֙1�rql�������-���#\������ ����խ���?jC'v��fB9Π�Y�h;�6yD�a��~?C6i0����#ͮu`ņOU�b+�����^��=�_�[,R[�f�13<�`pp��5~3�
�|��n��p/��r3��W�mSW876X'1:*��ݨ視�o�
��ƌ0'�m�6/��T#�c�5�����"�18mƻ�-��`i#�?g;�v��F�`d��Z��KVDV歌S܅'!�1!t9�V�ه��3	�fӡҤp~:�*�]b��Sk7,܂h��D���$.!���P|�n|��.\�)ĸ��͙�sLb��G�!}-���R�,���(ib���Y�V�r!JY��&9hst^'u˒K��$���غ���K���C�f��|U(`����]	o�Iv�T�@s�>V��*���x��/�pc�)e\��N��5Q�=T��������9w�C-!oߣ*Q�'TW�<�����������;>�f�<���j�Ȝ
�{�'��dU�PO�\}X+Bt���e��!�=4)�h5���-�?[M$�A�Ѝ���i���v�!`���)F+�"Q�p����.
��aU��<ּ�i�2�-�\u���Ӗ<&��d�O�'�T�PG*�a�hAڊ��ɘ{�C�U��,*W�¶A�K�LK�qLD(#����%�څ��� �q�ճ��%����ޑb}�{�3�F~�ၴ@���°p$'$��O�6�,�h#M}ꗞ�ʧ�
�l��ܔ�t˧5�X�MB���h4��v���	̘WL*��p�sh�(���6��҂����ALb~���<�L�c��w�$����*Y��g�6@���	���JdF̴�v����-ϳ����'�E$B2�����~[r�Uu�*�H<v�.o�f���t����2��:�N�aI��AUV������v%�W�����;w���	��d֌��f�7@Z���}��q��S:�S�'y��y�a�GF �>4p�hszL��c��������V�W��u�'z���]i�[z0Ի;�����>��X	3�"��~���o�)OKi�h8p�k
.��r�7��@����`�k�7m�gm��2ģ#�������:��{J���'8��iK+�?I8��U��2��(^�SsЃ�A�W�.J8;������[� A2�5cD���;���'�j�$�&�L�,R�/�X���&�b�y��X}Ҟ���j%���:���(f�%c�q"��ۑ�q�3h��*l�|qY�(����{<dh�F�8�@_g�P�C�#I��7��T矫g�a�L_.$?�q���4HmΆ �N�'>�\�[��}'��#�%#�Y���K
es�	�2�.
\RJ�*f<�V����u���@�
:{��-^Og~i��Q�%$W��:�%|M��: kEބ�B`���LACջ��IS4ܠ-oB�W*ؐ����@��9���}`��ы���Sc���n2ϗ��1]vݮ�޸��Ph���}�5�Q��[cĬ�r0eӵ����A�[�fN9���{��ƿ};<W.�̳�%�F1Pc�'�H�_}/B���fYr��ҁ�h��P�_��FV�;�YmJ9LK���ʩC���ء�A��چ6:><���Ϣ��;��*�g�ӿ��.��jg��(a��O5��}~�<)h�ψ����EO��؃~n#Ff��UM@?Ak/�B��=w�n�%>�#�!>��~6B��+(uU�ܗr�;�GV���|>�M������U�>�Z^�����.5�q�ѫ`i��P�ɭ��E���X�����L�R���3�.�d��Y} ����5á#�b,ðI��YG�L�˼}7��.&��S�u��_[�O�{� �Å	�ֹ�+o������y+��E3�W�U��AL^*����⹐��JVxcp)���R��ڧ�O��{+A�ԟ[��ǳ�L�x�p�.�(�)3�� �3���B�戎,�%�C�d΄��b�@�ͼ�e,�Ͻ��h�)$�
��w�*x��;Z�Q��.mnis�(���`EE�2T���9�U��N5u�~]%���_:jO|�(�� ��(�)o��@'6�}7m1�u�,�?��K��-;���� y����M+���b�?�b�8%Z̪3���>	�L�р�#�\�`r|��w����n[i֎ә��Y�U*G��;rƹ����6���\��z�V�>�M��&�����rj�����b+�S�� �w�h+n.�����3�P2��e�	�n���'�1��֝<�V��>L����F&��U䭖ǗA�YUb�Ѳ�M����🇿l�m@�:��6�É�\�_�d�u?�U01Жý���he�J��$��o�?�SJ�:�?� ����?	-u��M0#ˣ���MM���I�4:�,Gr���B\��}�s���.����|r�U�J�B����2d��1w��(��:$`�ҌmY��	0��.W<�A���znn�.9��y���Ջ?5gU���e��-���8[f��i�I�@bu�Uq���M�Wo���V�7�gz(6�M`�~�l��E�?��p����Ǳo(GР��9D�ɢ�ik͕��.֬�.e�f� ��da������b�:�w�����QVutGm{=�8C�au�C=�_��I�9����Y�[�8��<��*�L<0���ڍG�����ĺ��M_7�]<���H)�U�D
��e�kZ�
�S饍&�������j�y�l�\D!A+#8IӘ@'�Q��Җh�����(/@��;O��4ҭ���ѝ{r;�k��[�g�`���K�g܁�8���S�e���Ƚ��byYJ��
�%8.�4^d(Xitu��c��S(�CV���ED��(R\L;Y�����:�@�;-�6C�J愬���zC�TY�̤H�v�
�:��<;%�T�/�Rl����Y��v�sW��'%Sf��2l �e3��~~� Z�Y��O��S��$6e���*2����y~�TƐ���lro��r�Iҏ�!ʀ�>30ZTK>��p��դoF�L�r�ݢ35�a�+���Z=�i>�.� ��YVMLV�r��N$�l������V{"]�L9Z4K70��_�5�o��	��F�f��{o��c���PޫB�{8Ο�.��|�tޞǋވB{2d�$��� &rYՔ4�-�M�ea�lj)�#���Q���\�UĿd�s�����]���������-Vyg����vcտ�:c��TZNv#y-���ӹ0�g�Y��̓���Q��q�Q�I�mď)��M9,���t����	�:ym�&��%���Y}�JZ�UC�Xa�2I�%�ץ5������m�`I��q��/1zP���[j� �ו$�m�A�ˎ��Qh���Zv�Gq�<~�e��<�RZ$��'�@KN��k��3���X�!g��Kì%
�w��>���/a%`����J�쯄Q�&t��G�t�!<Y�M��M�|Ɩè!� �ݗ�t������]{�9���S� 	�mC�J�#�;��2x��:��v߁5���W����π`[�IX��;���3�?��o-Gq7�[*�H=A�{fU��޸x��i���Q�y!>�Y<j��0���$Efd�1ɻaޤ+_�ֲ�bȤ���d�Qٝ���%ek��f�����$]vb���ir'������؞w0���b�F�fC�_�$*������g���;<����r �Gɢ����"�y�'D�OK靣��uEe�߹�*��x�h��ә%L8��{vO�s�8�S���H�1�]��HwkD ��;�JZ>|S�Н讵��{Ҿ�U����Ո��c5L.z׃e�ao�i��� �b��{�5��ʍ�Q�3pf �ZJ~��B&�RC��9�ݢQ�:�>f�}��ppj���%Ӑg��)�dc�CNt����2����0V=���B�S�?S�|4�`G�?��?)xy���`)�U|�o��oى�0�}c��hU�Lpo�?S>�	�X`�-w�N��+���H�і�f�ߦOj6�=��aڴR�jj���E(���$nP�VaQ*x�f�Jf�_C`��-�����UW"*D��Ԏ���A��J"��;�?��0ib&{W�L������W��qzF����U��y�:���n*i�3?+�蘇zz����L?>y��FN�i-�~�G����Bb�t �]�!��/�Ɏ�zj�nޗ�ܴ<\?�^���n�`��5��4�9W���T eh���� �g�MB�Fh�H�����Pr
́��,���~_�t�S,@�$�<f�q�h3�Pi����o {�{���\�A�)�e�w-/�%��]L��ת�������!>m���Ļ[�;?[�t�):R��K��6N��?Mb�T\��y�{�Ԛ9dg���U�W0-{��S�g���LM�TMw!��Z�CnN�uI��%s��Z�!�Q�µQi"�[�?Hș4��n��D={������h5�"��T���uM���������e\���7�/#�"H�����~	%�z�@C��i�ҳ36e^�P8}����+�	Qb6>�9Q�L��D����/̑Z����f�'�kʶ�f�`�*)�7u ��p1�n!�P�PB�;��6���ܞ�y�\�z¬���Ơ'�v�3-)F1%�#�AqрO�rZ�"@l>?��Xw�5s���c$��V���ge���-˅�Gn�yA���`Z�� l9ց�����N� ��*|ݵ�g��	F�3�r������������wJʙ���������G��#*�eJ5'A5��1�NE}���/SI�@��EE�^I�|5��Ps��Zp���+�vl/.ҕP��&�B��d�p>�澠�;/&:6|� �[�(2�(S���/2�V�@���I��^���-�=����$��,�}b��k�_�	������*�jIĊ�ח�����{��E��g����H���U��L���X�Zn�9.��u�������|������A�ng��M�����'l��w�5��䛎�H�ޘ|0I
�x���E$���F��)$2�^�����#ȼ!j;0t �jFU/#���u�{E��(����)�ֲ�`@̨�
��գ�q��?nm��b3.���F��h���3�6�o)���pGg�"xa�AЖ��DX��2��,�k@�~iW�#�w�3�����E���:P���=�I�� ��w�x�_p������s�)K��i+$"TI�?;�粔�'�{�FW�}x�E�`M~��	������H�Y?+��2xO����J�t�	�7ו?���̷\�+Y���?��3�k�uإ����<��B��\��F�,>Z��\ =5=ԶY`�Z�{~SD����)d����/P�hc��G���::+@�N��s+@�W+]p,���<�^n�/9�a�_�\��mQ�5��dq[`���?6������y:tA��������Dq3p),����2���]�o�U`���=J�s@P-ҫQ������:�x-�Q���FGx͛�0e���s��Q��>~�"rA�lR��4H}�Y
�AȾ7�B�����o�,�U�7����fS��C��� 	���^����,��'�t �pϒAz�4W
�]\齷�s(�C��(����x�焍}��ɋ�%��,n�\#v����r`�9F��5?��"$a�=P1�yݥ��p%��,����T��/;��j&��U@~'�F�Oc��k2�1J ��� �����\v�c��i��<�f�P��X7}���.�	��#����ҧZ5�M�#��d�w�{�Qf����@�����-���<X�n�=�[f�T-�Y2�u,@�?�V�e����l'TTd�$�aEX���mIيv(�"�O�0��d�S��(4���4�Hgyh!90���_q8 �ޭU��Ǒ�T��T��5;D��!�^0+W�X���$��,�$B�����&�DTw��f>8}xҋF�G���z�����9���Wl�
��T��}��C;���I�D�$�6���@U�A$�;B���'ُ�X*�O1��+S0Q�Ѓ	��M\r�`�@f���<F{a���+�Ӯ��?����#�+bV�#r������ꊈn9���<�ܴؑPl��;��\sN'R*��=ӾX��L� ݸN�Ff�l�T��}�&3��D!�<x��&9���V�	����}�Ф�q#��N��π��:�O������r�`2�N#H�7��j�H��6������p䳎�YTg�@�o�`��c͇Jx���V1=�D��߲��/Ͳ}���Wcy>|_�d�6?#�T_s�>�\}�U4�&�Od�71��1ߥ�Р���yT�_��+��5��j"��I���X�D*��v�X9����9$~<��;�I1��}�-I��Ge�\��=���o�q.��^��9��ӥ6��?�ݸ�������n9>�a��a�h���J��T9xLr�d��D�*��W���	���>[W��S����%TA[�� ԥ���ДwR��6�_�V0�h�wu���99��#�л�����iM���M�I�Q8��,�J�<�n43���0㼤$+�u��+��OH8Z9���n�	_��>��DG��[�����un��˧�W�B�nM��Ð1'2L��f�)n�$ڿ�����a*�ژ�'$n�j�3�;b�"�L�Iֻs4&�����]�HL���qxdK;�-�����#%F�:�nP�ſ�3�l|�ު&��?e����ؗ������!W�0���=����Q���@~s0�[�4e�]U}Bcc�=�P��a�BM����<̴�2aV� �I�(�5� �������>�1U7���%�1Tln��.ef5�������l�Ǭj�a�����k;�\�t�?����ńe�y������vx�o��'p/4�V�S��u��K���-�v����[E��CN�kMWʋ݉u��uPI���f������V�B��L���C����,f�y�GqS$���J�|�Sl�'lB��n�C���p�x�qBZ���K�'�Jv6{�OV���T��X46'!
]��WvF���X��m���W@z����_�ƩonX3v�=���~�^���n��Ȭ9f�_�Z&� �*~=��(12�iPX|ᴙ�u��h�n8�����c�gn�i���p��4`L �i�\�~�9��Z?x�i��J�9چI���2�U6ɠ�o)������'��u��(��i������K0�[6���u�W�;��ʉ�TRJm5b4��ľ/y����&�W
��Ĭ5C��t���bV!�#,�-��|��UcKZm�!I�<L�i�NŘ�D<Ce�/^����A�˲n�8�C�T^�`�9�i�����104Φ.lƺ�� F<�%��#� =$�V!�F��)�����J�eo<�O��غg��K����kۆ��J���\qѲ�N{��o���ux���&�u�M�S�t$�-��ccݍ�������,�]�V�'S��)�۪�P�b�*e�$��\
�U�h���2���O���R��'��6~�Dvh����\�>�]�`��o
�������A�sUM%��I�X��U �%�y��%"��.X�?��wpV�H4�dڂ����,�a`2���ﴨPv���V�k����}��һ�u�_KڠS����@E� ����Ǧ�Z�	��h��{~��b���5������*]Ի5��t�D'P�[�z�c�'>7�W��#a�[/�����,9�m1� �s����.�sCK|��2\��IP�I�#�E5�1HB���;�<R���br��Tuo�䞧n��*��*�X����ZH̽�Uu�Ȋ�k�{�YO�����D�D�pE�����v�T�����:�MbX�[��7�����|��i)��`1,�����rN��kj�οN"�
3r��p�9і��,f��TRV��s��~_,f��=E�h]����_F~�j�}��4���lAff�~>YG����a�IA���aU{���6b��@�\�̼��|�{���g>�A>�["�e���P{5�>��r5R�x���vb�x�8��枟ED�N� �<k���R��,���0�E?�89�\�j��"�ڎ�Oj2���?��JI�v�����<��Q�L�C�
�+�F^�b�g�UbI���=��t��ڼ�����d����4�T�pT%�*"jǃ��WG��9���<���LsmF��n|�����;u.G[.��N� *fҜ
�����	i���6ĒS0��n>�]�!\�����%[���ggn����^�*M�:�K'�X���A��D�b%P`b�܆�ѺF�[�묑R$d�bU�5k��V���Ip}T���u�s3�����u4�C����b��&�r ݄s_��t� 5:4l�q��a�ʥ�f���ϑ%t�6kC����2��+��������� p�
��0��o�Ş�{�j�ጰ�b�7�
qQE��-��"��pn>y\�8։����/{*�����_F��g�2���"��q+���S�a�1l�b�)�Mb����nKu��������9Cl5TĖ�2�>{��H :�d�� E�����9ʞZ�2������X�>6)T�}����_Tq�y�r�����d�+I`8s3N���(K~B-��x�#*2���?OZ*��z�;A,g�|�s�o����������Q���J�� �*+fmH�LE�IV�9�������o����@����Ix��"o.iϚL`�Èe����Q��]0��ԙO2!��HSIȡ����${R��ύ��AaY�q)
o��$Y��7��*]����n��f?�ޘ9<���Z����7��rU�#���Vo�NG��w�����d���3>�j����,�8�L3*����1�-Y��	��]���[�e���eD5���������+�����gh�`����荎Ȑ��5���|\L̞g�MSC�+ `� �)�R�<�n5{�H�#m���u�M�=^t����J�ۂϩr�F[#��l�\ĳ�m��Cvig�B)a��M����X�
'C��-����5#/?�}hgm���#f)-�P����a��0"}��Y�Q��F��IĺJ�̠4�%~(m���|8�D6d��(b��>$ �;;)�P�]a͂i8[l[���>���,����$�1��Y�������$���(Q��"=�EyW�N�E���������g6��0f^�Z���Jk��J��� ��y�lJr��6�j���il�Y��i��Z��߲p� S��|S38��)�|>�!2�TWzE>'��Sp���bZ �j���H����������쐿#�;3P�nw���^P2��9V�q-���_���Ұ�;u�o�z�I(���9�gCudl�r?4�@s|����Bv`FO�}�C��p�s�K(�_u�0�r�x�)�_��t@H���*�@(3�3��N@��vf�[�mP�
(:�%��=������- �0�db�Z��@�/}|#��t�$�TF$�/��D��R�j�S����v���\7�!,'�9qh3d�H޶v����e\�8�&ф�s���@���h *h/��>-�e����~�q��Ε��+��֧��i�phE}���󥚽[r�h����h���.f=L�U�l��s��G/����#��r!����E��鉵y��b�%��B���yõ]�X�V���T��S�7��u���8.�IHp�GͲQmc��G�X.��ֱ{i�#�f��^���������?#r�����:�	���b�Ű��<AnπjĪ�J�Ԇ�k@��ojM+�����#f�f�L�G]8X��������fz1�4�e�f��$5�t����Tt�Tz��7])gϲ���`�\ǧ��Z�E.� 43	�eIU;g����I@WU�-��GTf}� 4����ww~���'��q�����^��Q�G��s���V���L?�*"�/=|�J@�n1'f������h�	�"RFm�L��}mP�=6Y�� v'Φ.�R�\^8z� �����ϖ���&5ї�j���<�`�"k�-�߅�8U�-������.5�7���K"��C�;��Hȱ�Nߊ��7�K{$l�L�0}M�,�m@7�m��XZ����\ᗃ㝶1����}X ��5�e����$��bۃ��k��kT����=��w��� }��ټ��Z�9��z�����u���A$���a٢Z�Q ֋��O��E�} �|��B	��QO�����IF=@���p!�VV52�:+��Y�%V�t��p	a��{�7@;�^ro�[���Ք�.{� "A=�)��'��}�Tpd�Gx�)�c�[���L~��"����V���Z&�\����|�W�wȤ"2��4#[�v�;��������	+�B�j,2TNټ�� ҁ�K �[ͬ8�m�֦� Q1"��3�8�01�x��%�\�����\PJF-	�1٢@���F�e���z@l7�7�4G��Ѽ~���ͩyv�h	`^A�X~��b��	/e�J����z*����TU?�	u׌�^����MeiB���"xx�<�l	p	��0���\�d�Oq�B;]���cTa�D0j���(Kt[-Y'����\A�E���o8�/z���	�Dh�.��/��S�|r��6����Ry�^W{�':�jO�]4�ʍ�7���ԸK�7o����c��4̶WQ�Sc��6�����V}�F.<�[�48J]��P0����C�1P �-� ��\�Ә��n�m�%H]t�t�����PdG�B�J�Z�J� �p.����CP��dX=�P?����8��U�p���9�B���3�^N5 �'$زx�FD����W;��=,�ʮ%�G�N3��.)XΨ^|�q�Pc�*�BTs\��;��݄G��C�SZ�䥰�O����?_����%^�
�}V�p�.��:!����n�;��3�`�gx��Y��v�d����F�&y$���]�\�����+u�`��<���$��G޳�s	�f��CP�D��;z��1�t �W�5�����9)u:���$B���0|c߳��^��~1}�g��7#���"�	8
�+ώ��$c��CZ���z^��4�z+zҡ�V�r�1��9��vD���<q�z>%V[mx0r�"ȥ���']e�9�@T�ke�v�|Y�I�CW�3[�ðkB.�D	�s��D� [��`7:�H��8��<�w���u��}�)�Adξw��d3Ħ����a"��!,QY�-�y8��H�=[�6��ˢR���O�R����ɀ��*lj�([�/�F?�� �C�N3��X��n��¬�?.GB�\���lf>?�����[bd7v���3���_�D������
�8�4p�ZK��� ��v9sx��EW:kܶe[�����L������A�8�c�t��;�L�v $R�@���z��P��s�`E��H���z��@`d�LY�Q%��=ҿ�����f�X�}��T\��A�
퇭��0;o�g��]��������c�í��h��n�b�ڛc��%f�ayPp�vh�KC�漛,.�i��ЦM�:@�C��Ŷ	li��4���B(����oT�X�wt�.�4]����6�sgе�Ϳ�� ��C�#.Z��m��)���ǽ-I�E�nN*J��N�q�J5Q�7����y�MY��P���yo��M-��,=�S�˒�TQk��N�i�@�of��$0a������8�ʔ�,�i�^S�{��8jWF/�!�Zlu6N�cSݨc<���돲��yo�:_|!/P��(�iYgЀY��ݬ��ٺ����r!�j���z�:�S:]��iT�K<�UJ���X��ɵ{��s�8r�Xr���E��\ȼ����ٵ\�o?�KV �����$��I�h�6�������X5�r�>� &���n�;��i�J���S�Ԓ����Ok�̐D`5	�iʦn\7�q�K�Q��Q	���^�<8�\��ozƌ?�a"����|�,��75'�s�\�&�3�\�m��J��i��p
�/�Ku�6��tr9_�,{��/U���(ָ��;h\�yf��,U�OHHTBw�O�9��Bad�7�M������R�8J�{R>���h�ǎ�tJ�S�`�兊��O�^���u������Ӱ��9�/`��N�P��ЖS��s���akQ�A��R���n۱$���^gQ�$���"�r3KQ_�ш�O�e��z� �A���S���dB��>�y�p�>�D�;��-��s��`�hf6�z���Ď��(�������ϡ�u�l�u;�&4�)�n\^�WA܁P����VnWA����F�H���[�(�޳�_���S�U~}���W\�D@Y{�,Q/@�y�B�>񘣶o��q6�/Y[\y���b.)���)���L,�6��d���Y:���R8P6���>�l~U[9.��aC���}6�q��� �5�bⰞ���P��Ѵ��::V�5�"��Ҋ"_ҷ�ة�S�X���G�eb��u�{l�t�3e�@��Ċ��&y�Z�50z�ݣ���k �q����F�:��rr�*��ޒ|Y�P�g��yq���B"Z�R1q�r��4"��/�+�O6��,x6��8L�G�Z#�u+n'�m(#׊�Љ�68�G���B$פ�o���XN9��\%���*�`y{���#㴘�ƈ�F�:�<G���R���"���.9����q�c�����B���h���\g�{����J��(C�Q9λ�r3���PCa�����I\X�׋�%��p/5X�tH���x��p�]K�"ԍD�2p����f�e�{�"a�_�%��.(.�~n,�~�@����Uzw���3�k_������n�A3&�I��i�ʂhV 4Vső�siꕫ�2�QkQ�&���Ų�%,����i��M�^kk($ǲ�k�g�!�%�@5�= �Z2�]�܃:�Ӥ���B�pU��R�\m�e��F!�2C�%�J2<���Վ��ͩҷ�X�J�~~�c�䟮ݽ�TQr���r��\�Fyc�:��Ʒ^�K/�R0��{wW2��]^��$�.�H@����%i%Sh��.������B�׌�~�ss�7�45�wɫ+�#���5��/9�%�>��!�)�\}7�����eb�D����L��;yj)�(�g��p[��ʓᒧl~�@e�}B]��3$
�g��6]�-�d�9e�C��U��̳qU��FeC���8q ���T7f6F���?s	a��ς�&��g��
�4O���	�^��(|����V`g�1�V��f�ࡖo�ĥ���+�Mǚ��C����QgTn$G��$�z(���FK��Nin�/�X7�?Y3	�4H�w �W!<�r!��Xb"�C�k�����c;�ݭ煿��J��� '��j�h;2����[���@�(D-h�K}�`��a8ʧ�q&�׍yO�F�Q%��M;�,�1a�/X���Ce�����yp���^C��U]"��Fn�Mڟj3I��Wy�}�'��<*���9� %�T�ޜq��ޱ�@N4vtIrW����U�f�L/�Nq�"��V TP6ڌ�������vj*��*/{�aX�N�RH{��B��K�<����{ܠ�:���ᣲYh��		7�9���\2�9b�G���Z�m"�x�Fh}�7v�F����x�U�����(
�֜��{���������f5�+pP)q�R��n�k-xT�On���X�dg�@o��
6�W� ��PO���[IiU73���m0�%��UP?�&�#�Kz����]ֆwk7AY�\s�i��pS%m�p�;�n�`V�HQ|R-5X�YY��˨�f�����+Ȋ����-k�,���:�>�����K�rm�sԀ�|0�ڐ���OZ�&�4�o�CG"?�jh���}GՅ(�T�M5�hI���%a2��붜�����r�0���`?�M��2V: ������3�H+���F�@��Z���}__�|A}ډ�;��O$��Ln��������Ue!5��2E���y�7ի�W [!)C�M��|$��鐩�g� [I�����D���Ԏ��[�.���"F"f�����=g�Vٝ�[+�u{��
 Z
xA��Zj	5ŉ�+(Ӈd�?��cӱ+n��GObg���<�i�e�ǂ	׏�	~��5�U=��	0���
i��PJ��?�]b�>!��^J=�*�T$�zf�EeHN0��k�+��pq糲���4�iz{���}�k�`	�O��N�,�q�:����؃1h�!���8Cθ"�j���y�Aԣ�f�~E�=��]?}E���5�� 	��;@7�gt�����[Y6A��,�M��l�K��e2/�_�6��	
�$�p͔?������9�\����L�m��c̶���d�G��+�}q�Q��K���1�>ņ�~��+��I��*t[oE|�)h�Fڋ��K�C9�K��Q�
�����U�H
9���,�'�e�\{��"��Ach;=Ѳ��M��Ub�P،Ԭ�j�3�v271\FR���葀���<^~7%	�����k��q3�l��W�	=r�ȗ�3��ئ�{�q�����A}�&��]`h��:��p��B.T
A�|�y����.V�o���.?v�?�VD��NK������ڡ��W�~��n�@�ذ8e�ԍ��B��=l]>�?�߯�6.�\�`���y��9bpC�~�9b~	��������uL�4��B����9��O>�f���)S{4dJ�$.��v��B����y
LX�Np_ʄG��<�!��LQk�vb�2��O�A�����"��IZ^^v���=�1�1�|���eY�d���g0'�S;DΡ�0���b�N.�+�H�_������t��	5M�BY��j��>徥Ύ���?��N��P��Y"	����?�S�Dk.o� v���h�*��Q��\�/`"�Y����߶P��,$����o��a�T}�����
��/F�S�my�@���bV~�����}�;L
����6�C_�p�?vE�'��~>3�@y5�����!�wf���+�y��+ ,�\]%.���W^�v>�o�R��K�W��ig�r�L���3/�޴�����̗y��։Ek*���^o�q�l��LFO�
�˅*2l�=��`& �@���;�5�˹�wu�T�������w�T���f $7'+�q��{gJ�aê�I�v�t��n�
�@���ԝ��	,�c5)�'UC�3CEY\��
v6�!w�)릸��V̢��B�_��j��b��t�z^bg9eX���5�V�T�V���>�<��=�}��W�].�^щgQ���4�,u=�4)�7��-��
�(���U7$.J��'�lv���Vv9W�,6�Z=f�ơ���X]��J��γ9$�)�37�Q�c.�ь}@��d{��F)��j ��?&�ro���@�N���FA_�7'��sy�<��.����2�����N �G_������v S;p>���zx��/PØe��L�i�0��`*�A��z�`�f=T�`�*ݥ�%�\#��l��F�`!��?	���2��UK�8t�.YA��q;�\)�ܲ�2VN9$	Eͽ�}�P\���T#�=���+�U��*���F[U�Q�s�'�_W���ؾ���;����j�?~ѝ�gg�\�4�n7����ڏ82�jGm<qW7��畟��QN�d�3��R�u)ک�,��v�	#�6��xn��+��2����w8��?������ёĲ7��/�/��{\����]V��"�a9���z͸��ģNc�ܟ�ގ������)i��N�:x��`mBk�Q7j�1�j
��s�?���#1�|�/�I�;P��4YY�X�&�H}>�馸�{�cPDm�VF�~���QgvcP!ĝC��:x���t3\�65�����������b��>r������W�/0PK��17���p!��b;R�@�z����,�����G�����Z�&�)z�-�C�0�ѮU�~���B��E�т�8~����73C�μޤ��7�#�ѫiӋ�c��N�I�KdZ��M�}�b�[T@��Z���,�"H<3�2������{�i�%�תCm���P5���N	��J�
n1.�LRh�p�Xv���5]I.�������><6b*�80��++�QP�	������
s7xS/z��*�q��2:3Km����mrhY�I(P=�5��1΁�+C���C��������y�%{� "~��l�[����sV�U�%�X��uU�0x	~�n�~`^�Y��\��@ڥ	C�)8�
���t���sc�v�-�r��`��:,g´��*��e%�ޅc�(�gԀ�l�h�fW�a��J&Ր����=�B!i�w��"��50=%j�%��\cܤC�T�8^,���k���$8�mA�cѫ�Q��gv�<��Ȑ_�H�h���T]�/�	��kP�(%�]`�JD�1H�N���G[G+�W�X`�X��&��x����P(��v�=mk��FtQ-o���DY��kMc���"qj��w[v�8��0�, �ܧ�����7�D��M+�S~�A�w��+�����C��B� ��I�1y�������i�v�!�=Ա��V�R�5pGª�r�=+�R5��;a�D��j	g�\���ݡ'��zi��'��:����^�e�bm��p`
�T��;�0�e���~?�G�a-��ܦ�/w<w�L�����bM)��n�	��[�vBJI<���׆}�)�"ò_aw��N��p��V�v�J�F;�)�ԟ~xkF�����asHz&d־1L�QtO'�ܞϱ�28�A'���I����ǒ�z�\��������I=�փ���[���J"kl��Eh��0��B����^�O��ԑ����F�N�s@ So~W�a!)�g��	��8#�8-k�S,�WĘȠp􎅸�K�	�̚<rx�o��m}i����O��&�u��4~4�)r��Ӏ�"�,�pB��R~�a�����_����������A� �3	�����y���l�x\�A��_8�[X���1k�:�pգG\Hj1A�J�і{�QGX�jj��߷��jtS%��֓���& �	]����o�v��vS�+)^�s<��l�A�)7$����ϋ(ew���Y�|�5�5קN���p��� xI����I�?ý�n�[v@�,P,j;��j6�T�*�Q���o�^�>+�"�cI�ò��Ѵ\~Ȑ,h�Ze�_W��aYs�3/1��ߺߜ����1q��x�;�Q��*L�O+"� �j�,;���ђu`����L�"�����ѝ��������B�K�[�3�.��Q���:/���!�Aw�i9�/j���:�Zg&��m�CMo ߯ ����ć�
�uۦY͑+�Q��N�#�
���r�W0��7%;b���G��f�)�@)����>Jl�/_�L�L��Ĩ�5�k'q��T�j�1�9:�2�̌��h�&�
@7�^�*�׎��C*���m7$M�c�WA�o��y�������� ��w\?|vڀ��}�<�:��F|����u؈��Uo����u i4��v�*��l<~�߭F�����9=������)eUцU0�s����A�|�ЗHVu2t!7��	��&��[��3�,4�h��d�K��ɳQM[.EE� i_��A����fCv�;��q��Uu�G}טf�Ô���I�!��B��H�j�d�Q9Y�*Kq?�2ٞ���ݶ�Ӓ7�RH1��+����n���e�@ '���uZݕ�}�~�=�H�,Hl_� ��녯4	��EK�<��I�&Syl���ju	L�9��1��|��P�z/��X#>h^�
�oG�W�%�)�̇F�+F�Hu��[�p�I�Su ;��&:~l�w]�$�%j��C�����ع�FAo9�3�V�d)�ǵv��\Y2���hɴ!*��/�?y��B�+rp��2��x�{��o�D�z�āv�͎�ѯ�p��F2�I6�&�/?�JꛦX�'�wԪu-�4V�0�/�ݒb&!��*m:1�L�9���*)�Kb�wp�ր��C��Q�lL)#X��w6w��ä�-��u�F�D�hZY\�A�t������w�a��q�T��{�}޼inI��$������7���ls�-��}�ƃE��odF1S?|.��lwAy��F+�Lt?g?)J�:Ŷ�O�����7w�6V�:�9T[�
�.:��]ƭ��y�H�:�L����㉄$����1�f��'#:$�X�j����_���DN\����P�N����*����r C	z��4}1i����]� ϊ����o���$�Q(�6b��ˋ�E Ѥu;+� `ӏ26u�����jB��0\�u@��w��1��lBAOk	F�����Jd�����$X֔J�u��;1��|�|F�+�;���vjL�$�P����+'�e`{�߫{ý.��W:.�js*��:rMˣvh�d�z�u/	�%�����E�A%�ܾ�M"A�E��#������J���:`���9��E��[d�h�^�P#��)ś��Ѝ/J(	"�_����K2f�mtP����f2��W���wXDh~P���V	G��z��љPR&��epb̰�!��\?S���X�8$��Yy�1F:�+��A�O����Pykx���1'�(;A�?�}#�?��T��Y.�*���C�P��������)��Hu@�>8�+(���%��� V�u����겹� �)���u�5�S/�*/��F�T�z���2��g��k����_=0���U���R`�<ˢ�19ދ���@� ��h�>�3c!�j���tp���8�6��:P	���]\O�a|�b~ڃ�*{����ҭ�ƧC4�N�B]�U� >�8��s�"�E(�| 9oD6�6B��k�d���
���l�JD��)��"���7ݫ��H'�KՊZhQ,2���7\ƻ�v��";�Č�K<T	^�sK&��p�����5�g�!��L���������K��?=��2�Ѻ�ߍjZ�UZ���|#�&��	������,����&��p�������-�g=uZ��E����xkZ���K��K��7@j�l�Oȏ/��L����YH�&�z�����h���(����I�_^-3Ea�͹��P��7�:��;D�e�~[�]����z�]�I]�9�	=�X��G{�l���+�\;a�o�n�֡�;�a���g�������H��`���-MgK�t����������[�G�med|�͑�:�k+㵧구8�o	�@�<t=�����v���.�}��������t��������p��I���
Z�F�d���
2��v�M��Ͱ,3W��o���F�&����'�K.�'�H�PL��&�ăRC��}��ѐE��f���msqϦ���VB�mn��o��"c�K'I��Dk&|ި���tci^' ���sB�(��i� (
���@(^s��~w,�����d��W��b���v�	<P�z�MP�qZ6�4�X��_}��Db���!9�1�U�(�[a������+��Zt��h錚�+c`3��k>������s %Χ5�rW��#�>���~�aՈ!%��	�y:�f,��t9��O��Y�w�zI>-ǒ���-����O�J���+F�@� �.ԹqO��1m �Je��<��A��^-h��!���K�]	�u���0UN�}�}rqoya���r���%;C��f1;�h�L�Om���nɴ/�@�6�cGWl|��w9�`�Z���F����9/���4����Є����\"��vt�0�����v:� �ZJvV�tU5��!��!!=�s����+R~˚�sƓ��)F�7�J�W
�z�?��x�;��B6���"�l��2��/Y����!�EW�3�TDֹ�<\n"�-�.�|�fk��P�]�m������f�sH��XA g�q,Nj�ub���6�@Ji�0҇7¥�F����&8g��U��!#�A�3�&�3�E<BF�G~��!Da
"���4p떂��*�rh*�2�_��������u�(�e��(�� �|	�]<<T��`�#��EBO�z0��ީl�^&A�S[���n!U�	��	2��'�����>S������񶏐��d�Ct�=��º�p�B1�#�[�}�M���
����S:1ˑ��`0㫜Iإ�\mǋ��3��Q{Qc���qy
�͢4����v"ݜ�P3SS��1�+��$n��wD��ľ�[\��odB���-Ƀ0OXz�zۃq;P�z�E��!G�<��#p�975�H�ӻ�ܝ��,�ᑵ�ws%�)Z0Ӿ�N���^��* ����41��t�(��w�*�f��//����#%���d�u����
w���Y�����H{�Mu=�g�A��YµeѶ��c.�-~.u�vK���	����4n�BݧS�fuT��#.Z�4��YFr/��Hd���0@M�J�!Mժ�p9�����i2.N_��F۱����/|v���U���t����[�1�4O���^>�X�^�@)�цC\T5�b�L�h�2��/Y&��3�تlG*�q�cJѼ��ԝqw8�fK.X&����3'j�Z]�w���z�]��:���30���C���Fv��$��¬V-7�5s���h�x�͍�o�����X���3'���q��Y��l�M<5d��u>�p�׎�[)�l�W����M�Tg&����������VeV]`{�Q��;���׀�X#Hnv�Qd&&;]
X"*����K>�r��F���<�dd���n'K�FCuo�`��=��!��-F�����@�F?ݺ*0s�?6jĢ�6|q��Ɯ�vj�%���pb�y��{0EgKP� ����L�T*�=��g�M��	؃IpOѤL��z�"�l�[�nJd�_�'*W:!T��d��R��Np�.i6��mǱG�VC)�,��G4����p�SGE�s*%{�^0 h��*�RF��ޠ��y�c�����J>d�'ߦ���L �Ep��	*�< �sv���1�i�<����q�[j+lL��t����j+�?>��i �S�B���6�6U�Θ;sV�˩\����l�`��;��餕�+c�Ŗ���`�0���#�i}�l9v�����-q&/L���g�dl��Y�d�}W�8��1�+
NѼ�kU ��/�����j�ˢ9 B����pw�d�a���!���S��n���z�Wk��Ĭ��.�� ���}#��,�f�z�22�͘���T��	:���$\Lc'��j�aZ``�x��cS�q�;��~Uk��
�̰-���OD��J�I��r'Q#�Y��7�qlnoǬ�qN��Z,kp>sNL��S+��@m��A��c*����j�~���>I��g�"���q>�)<�_:y�~l2��[�cH���AIRT���`�t`e�N.�񗒘`~X��=�R�Ys���-�A�%ovW�?h(|��:�Xޜ�_1B�J�p��g�<xo1��a����5�c��NK
�}�O'���
q���u��*]�9�=Q��b(`旲]\Zo��ō�o�F����&Ta�1�b������k��]n�����Iiξ�<��+(_ߛ�_���ۿ
�2�}KRKH NJ�}��3?�tр�q"U��r`��l���xD��;�Ԣ��{�yM�K��9yN9W��a �����r(g�>���_l|խV�@z���FV�&X�W��%�����ˢ���!Vb�����a�D�*�'���F���C�8��7<O]�VߒW#k��m��]��&���!jND/,�d=��(L������mU�oɪew�R;�LyH���n0R��!���-���+/������Fl��=��"Ζ�3�,���G���`w�(���e;��Fe^���5�����AT�m�"v��Ⲣp����>����ظ�#���@q�̎�j�ҩs���_��z��7QRJ����dB��J-W���S�Y���9[6�a:G�c
���h�D�A����-ƐT��i=�U��L^VJ�m|NfZ�.�:h��)�/�p�`�:G�J��ǽ:D+��+�ᝏ�*S;�Pԛ�jp�JN)��Mr�.����6�I�(_4h��A�O�s��-�S�s
n�G^�m�L039��sNn���N�H�̎/zc���h��~���7�hS�l>s���I���o���L�'n*"EE5�H�W�4��!�xa9ބ�N��C<�x��!6a�����Nz�C㧆�%+įk��<�@Z$6�/�&zkKm��~��ӷȻn�EY��0~�qψ�6�#��1~A�#�n`wB�Xx ����#������7
M>s�Q}��F�ٟؔ�D*Pd'����L��3�D�҈X��+94x1L�X,e�ï���
�kJc���v~5��Q�S��Wo0�,�[t*|�<�-ٲ���c9#�=\& �Sa��lQ�ynT�%i��x3���#�sT���~|˒�%r���B(H��V���=%���ImȒ�Y�^�����բEL ���D���,�"s˯c���ɲ�HPƐ�|J�߃%��?�:x"|��C���Yc;�ȇ;~��%�	�;��U��HO�l��a��>ҁ"����;d|�z�7m@�g^�N�kĞ�_�Z]��^�Oį���sP�ǽJ�i���GIK��Z�"��vևh����੬n2�we"=�'�y�Y�6E0�Pmq�T켜�"�w���/_��1��wDA�x@�Yr������oZ�Rj�L�`c��I�ز����df��#Q!��ߣ	�8p`6U��<��ð�� &��>[tqJ���wH����� �]��*vc�9Ȝ����q3r���k��©g%�)&���χf�-�iQ$���܆�7�@7-V��N�ko����N����N���N#[�}{�����V����w�Z|?��y��Xݟ�W�*�:FO��Awr3�����ò�� ���9����	�^�h���`�o�G%���So©:XnHڙ:㥔_Mw1!���K��e"�"۬fH_�x������D�&Ò�7�a��#�h�3�8�2����5S�n/�p)k �V��Tx��~H��{p�,Qc��9½�0�­��؞��Ȧ�'�I�v��Z1��N�������"�,���B��@���	�?K�)lSGd�,��˼�  G�X�H��H�3ذ�ѿֶ� ��%I��p6.'��DҾ����w�fF ���vQ�T���F�I�ڐb���>�	gP��m!é8����RV�#$�
S:���2�|�r�Ve�I��5�	��&�� �O�����(4>��T3�wտK��}bR))�H�4WI��b�#vB���L�f���h��ڟ%8�K���q��*�_���!�?kIWn���-9SJ�/	p:TJ`�n׿E��zm����λ]�S�UFG����@&W�,�����x,��Jb&D�`}*!ijr ,t��%"R�"�I&�׾�V��`�t���_M#�?yt/ǀvQ�~�[ؑ�6��\hQ�Eab�x�m�T�(�$��+�YV�k)�3�N��h�V�4T��\�5G���Ɵ+Se�R��r�'6(�hQ�1����~)I������ۤ�A�y�gF$�&ض:Kp�)�@u�WF����Lh�,��L
MK@_px�d���ne����H��e9*�S�T�X��D�W0K�C��� ~T���Ǘ(tv0��*p<; s/�	�NG��C�K�J],q:�t�Q��լ'��v���-�"���ߢ�R�����f㩺������C�fǔ�s�NW����Cj�[ڻN�0��HWG��y��riM�]˲.Q�S��Q�Y�$3X����.��'@�P��K�M9�0
�2�Z�C�>��"8%-�Α���[���8'h����ɲO�f�dhT�s8�l��!ѕ��V��˶��g�U�պ�%�9��K��j��(x���!�Ȅ�L�A�!��1�p���ڛ���^
io�ܺr��F�!��D����g^�\&ZPP���I��v')<"T�;��O�s�R����k/��w�Y�$f�v�����P�{��fa��>Sm�˔�,���*Jj��)���_�'���)�wT�p���4�+ s[_�*9�чާ�-��l�sΕ�\������4}1��*f�ԅE�#_��	�5c@�t3�j\D:�ս�9P�k`�*��(��u�A�ǥ�X��8OF��'8���/]w��S�3#�ҁ�5���>�
��j���Q��p>tj��g���[�QS��{%�g�9�yZi��+ܙ-�R�zޙuZvBq Z4��%հ���E�k�;����R��XpH����Z_�-�#J�h�\�/����*��x�x��>��8+�9�N^�7�m�f���l$O�L,y��EσaH��pNN}�mOǹ�1&�눇�C��B@M֦ڟ&�	�c�<�[l@O����L� ������ӱk��X�j�Os����OԚ2v�rY�RT�bE3������� +b�:&O����
8�w� '���x���=�M��Q�:'_��,\A������o�tBX[Ue!?���W���*3��w�t�r�2���T�������t.���Ih���'�D��5AV�˼�>R���T��=�T���.<Eޖ5�b�-����"��Xb4�^�ZkK:_!�ס���=�
��d������3�^�:y���Z�ؒW$�1e��9Bn��6P1[R�yb���Oz�[��}��0i9�d��5��^�tl��J>�y�ə(!#1�����O<�װx��t�0�E��u�Ņ���[;%�a�:B���K!��K2Z|�����ReJ��4�~���*�\�ҙþ{Ii�Bi}���r���V��#Eޱ�1S�4{b��R��
O�@-̈S�a}#D=�?��Qj�3�Ǩ�a��<C�1�� �O#�]���h��(鐫#��\���Q�M/�jiJWI���6N	�	'o��W<I������
/�X�� � �AM�Uț���R	fJ[p1��Ծ���Ra5��w�3!]PA��Bs�AԳ���Q�I�~��ryT�W�K(z08������+ގV}���.f�v5Z,$_�1v���!���wSr�Е'�b���0�*��FE�	B������;��ͬb�U��O�o1|j���ؐ�-u��O5�u�����j����W� ���NO�"N�oO$. �830*o��7�&v���"�ܽ:uq��e؛��y��"'��˥��� ��ȓ�va���Fv�o���Sy9m�m���:T�۽��`�X��؈c@�i�8zËX:Vݱ�c��5k��빕2Eyv��v,e�d3�<t�/_�f��1��v����в��u�H�	��H�=��C[6�*T*7�K��2C�d�!>�H��|�=�X�>fqq*���li)��2�W�!I��dE4m�������ۭ��9�!�=���D�/�G�>c�D���P�F��f���T9+�pl��}�Ke'��w��?T��1�]�t ��֭O~���M߸�#^Ȱ/�.ch{p��J�R�Nꯦ�0��[g1O Uu��l�	˾��L���fh�g>zNU43Y�:�w<ΦRӧ4���,5��x�.��$8��р�2���T-jc_M��Dj>T�>6B��!��S�&�8>k�+��X󡖏��O�6q��v9G��&yZ�Z7Ho=3���T�O]�ƭ�^f	.q���Ey�7mU����l.�m��6K�#|>��%5����N��(IÃ���>��_��l��6����26�z4s�#4��I�!M�w�䯴qV�S�S
�:�Q���T{�uK�������R�$U3'�/y~?p��K�.od�4�J��a�ҵ�CF�,A��G��e���v#D���(����ڻu��%��zOѕގ�I
�N���H|h���-���"�4�p69��I���ֳ��\�1)27�A�v`�fW�������&���
!�m^���cvO�Gv@������@�'/x{��F�ʘv�O�s�VS�9��S�~�>`^E4͛����9IV9��д����d�=`qM�%l��|��U4�#���(u֥%�_nc��<�K���UA�)%��M퍁v�|�ېP��r���HAۃ2�tS�\����/�m�ĒLb��Ľ݁	��ηm�=�;ω��]�Q�J����!�*n@nשq)ب�E��Sm7����B-�	�E�X]o/�v)���k���L�j�.}��d�i�Np�
Ǽlħ��E�&{��D5�@�~����~�$�:+��:	s��7�9�.��x�ĕ�C}�&������� �~f�緅�6���,G�<Wk;��J��)��&��=O�g3gX�CJ�t�rm����?(��,C���p2;�ف��|�a����-[��5�x(��?�E�#IS:�)�x�κt�4�����ƟM�W�G3��aEF�N�|8-�>�߰L�3�:�|(i�hL8�����;��yq/��J�0�.҃�.c]�R���c��:��6���Q�����-�ul�!��NѼA�lHN>)�4���g�����[��dķ̶��^lm�{�a��L��?��b���<��;�OWکz k��
]ɆI
�j�Bd%���0	��<��߽��G�dE�,����n�:}�.:�q��h�|���X�af�\_�ɘ�|l(!g'�? =~i�a��L�����<�� u�x��E����]&I��?.zw�NY��Ua����V�g�m\�!�^�J�݀f-�	���[��I�&g�&���׻N!z�v��P[����gę
��y��nq5��)��&	Sɖ�lӶ��f��T�O}���������I��3k�%#O���M��6G�Eܛ,,ׯv]
gy��<�J������)�F��D�G��
ih ͊-(/C��,��H�v]-�za	XHS�Z9A���øS�T桨G n����h����K�}<����R�Ą�b�".��c�	��A׿�D
�e���ĥ��S:;��:W��G�����9���l�լ� �~F�+���%����M9۳��:ծ� A/�86l[��Pr�.����'3�r 8�1�<��ߖ;N�%� &R	�2�'M�z�����\߱N{��I&�͋ێ4z�_##��UV����HR��Ҳ��}fA��J�@q�I�o�u���N����6��8!�/��=�sR�^��Qf�&0���fP H�S~1�)~��sk�.��H^������8��ī�e7����T��`�����t�?V�!���W����q�`Ώ_�j��
ln�W��^*-�s�В��n����-��hf�/e�����[n�ȹ��M�4�\�#����(@d2X`�K�0}dvB�����Z��+�U?Y�U����ﳺ�5�����H*?v����&N��}Q�����ʊ���4s@�1�0��$��#�,G�'?0��.v�2a��ۀ9x�ͼ�{AP���I���[}h���.#�}͚q��t2�T��*��i�!A���788"��8�+��q��r3m�A��B���MщT�,ueA����8n@=�6/�M���Iu���X#3�S�ϸ;`*��9����
t�?s��+q�B�R�O]�sl~y�]lL)N���-�{:�s��_j���2?�ܭ	m9O/	�n>�5'0l
&�v�w��ڂ�(>�==t��>��`����lb�dt�?�'��T�ʏ�^{n%l���4K�����sb�1�Et�Mj���Bt|{��nk�j��H�j˟���A)�ޤ���r`���p�Y�������R:�'E5��#d���deH�wo�Ӈ5E^���	�>���YH�C]��E�j��`SF?��^�i��ѓ^�Au�n"ZK#����XfBMW��[�l�����Pq91�Uź&h��v,���JCs?��2����Iߛ3�.����o���Fy�y�/�.`A��!x��V���i���5�yW���;���s�P��������q�#F����(K�Ayk�o�7*Վ����r��7��5g��1Gf� j�pK�t�.K�Z��`N����H��F��mt��?V�: ��D+I���y��d��:��BF�� ���q[����c]�Z��R�?�kRb������7&�M�����T��W�f���|���s��
���U�t|�0����Y�bIo���? ���
LP�)�B���	-�A����2&�B�.s�ǁ���� ���)u�\�P%z3I�遛]>t��HS�~v���Om|�cG���9 B
���o���~��<|�}�s��D�1�m�\7���$I��L_���c�¿��<S�S��M`���2�E`�Fv��x��qF7�Q�9i��P��㙅�9��/P���W"��^�n0�b�nNs��4��тF����>�����ng,q!Q����ܦs)��${p�63"��zK��6�,��zdc�:�2\�������ϊH)67?P�����pj��8��ƞ��TV!A��U5���Y$e�~gKwJ1S��bO>^E�;��T�Te.��^�,xTT�<���Ԧ�t<��-x����/�U�P!�_����|�ʏ�g�OM_�h����*� Eo��N1�����@��ۗk?ޏi�8�"͛��uft�M�TX<Ҿu�j�������	�7��~F�>�<�aM|v����6{t��;�Y�2���N<��t�x%�ɇX˻ژ��Z�	�L������ҸOCݚ�(��NB�M 8�c=�O�]j�[w�e���j*��9O��qY�U�%���#����!G!+e�
w�=�ι�ϳ:gt=(�
<�]yh8˳slE�Y�A%�k�%?��G�����R�x:�&�e���MqTM�B�7�:iZe���5�5�gl� �tC{!�$������(t
�PQV N���C�u;ɾ�ܞz���}��	n5yY�C��p��B�Rف�tʌ	S׭�2��F#���%���vy��[n�������n�uN�;�NU��;�c�$����w��j��$�Ƌ�`�-5�P)��4F^6���b�K��E�|�=%b����@���{��x<h�窴[�6P����ӛ}�[����XG��� P�+v�N=�s�öQH;x��'�ͱu�,���F-ѥ������j"@C�ą�	��r�8I\���j�Ut�G���J�ҐP���$�(�i��ax�-���h����gW]�U�B��vD`x�F$�VT_ηr�I��ҡ�A�I�2%ڼn.�zӹ@��*��\�Ǜ��b���8N#|flCG0�p~��j�^���-E�[)�;�J>��G � ������7�>�Cj̣A�T�o�:��K��+�ts���&ڇY4=h���!���k����}�ʨ^�[<��F���G�_0rN��9kz�.o�����3Q�R0�T1{w�����&ؓ��R+���Pa=<s2⪀�"��'�'/���kW�W D���Q��jK+&4M����5"��9���`wˬ4����$�I��X9W��8�I��M��QRj��I�� Ӈ�Ǌ+B���آ�%"#NK&���ɄƇ9�k�ڀ�}�Ҍ��#R���=���Pn��i�2�r�PA
IHq{�<P�@�V��CBAs/�Uk�PQOd�/^,!��y���;ž�������6_PGDe$����Hi���Ѕ�.1|�������Z j.&T����w�g�II�?�N8�Wp0�0�p����!�*R���<0�Q����ڵ�V+3ԙ����������}+����1����w�8��8Q�܆C�o���,�8a���{;�� ��(#�.(����k �3��0M<���w��0؟zʻ����чkʀ�0���3%H��~A����=��
��g�����
���n�M��*4�}SW8��e(��P�'���5I�̥���ow���B*���\�sq���l�N�����i�H���n�BQ�-=$t�7�}�m'��2�q+�� S�[�fA>��?��æ���"���<^3���7eެ�]����=����2�V�vG��{Q�D�M���9�r�a#I#ځR��0ۋ�'H"m �i�Q��1Ғ�<��Y�݋"NӇ Z�7����J�Wy���
Ʉ�
s��������X� ^����'��"�U����,���y���[r(B���&I�g���"@Q)��G��;�$��l��	����9{�`��2�j�.��<ߵ��d�;B�<&����ya���@b�>�6ƣ�a9�'��xk(,�#���#�/�	�J6�;J�Tt�ؐ�ޞH�P���4�[ܽO'v���u�`1{�L�u;lE{�b7��	�es!A�{!8�@��2+p��c�����%z2�_��h���\`Em	)�ȝ�t�045(9UȻ8Vآk^��iV�^y�����s�u;�4�b�v�;�V�ix�/V6��\��?�	7����"�v#���[�=C�C�G\���jΜ0�PX���>�}��ό�Oݐ�mˡ�fBn������Fq��I,U�PKe�cm�f�D;AӑuAq���xDe�Hҏy��H����刜��(��U�{�6h���rG��ǪM�<�Al�3���s�(��rN.���T��{)�y:*����@�m[�m�F�t�)����ЗM��4�����Qx++��񯟭�'��2�|�S�_��mj�=Uei�M� 8��,����o��H���5V��)ܶ��}g�YRU���:�A�S=����C�|�#���g߉�m�����7�ʮV!5�EiMg�~�]o��1Uҧ�����6��={���M�8�9��4A!�oPG�(��]q��2�S|����'Y2��A�I>M��mw��������덓]��O����ʾ�n�4J{��o�lqW-���i�ж�2z��^KӔ�~5Rh�P���6F��8*fֳ�w%.�F�i�?IuJ5�����������"��gۄ+N-��"���
��?�9d�zrj�lI����?�S�5�tcː$�\�+hf>,�Zf�"f��_p�6����i��g.V�L���t�b�(���5��0ZFP�@��/���<�l����2>t�����m��i�����Z<Ok���\	����Ʋ%ǿ����^���GZq�S��H����c��`&t��5��Bم���m;)��:4٦i-�J=���_gX�Ȫ�]�$��&�e5Tx��;O]�]�܃�a0B��Q��[�9Z���yF` �hV����T�K�8FϿ���sm]���3�c���eK���l7s��\Rku@S
����~Z�tRߓ���4���
m�7���)p�~����NU�n4)����^�Mx�)��xB5 W��W����\x���ϵ��$8-�51&$E'/���P���(� ��ټ����ߪp�iԧ��j �Vܙ�H���X9������Q�={}r.E�W���x~s�jD�
N����I"Ы��[PH��,�]�d�F߽��;(	_�C}�Y�u�(@vNh4���Nx�L�m��e�G-�"�z�y 
&*�g���(�!ezm�H�_��A'j�\�@Dc�|�K��/���T�nÿD曡
��e<�l��� �몐��}���Y�B�g��	K�ʅ\zz���o�0e|k����!V_��4T.{u�P4]�n���]��!�5�;C�a�Y�*�;�	�fF֚X �}��:�����2�_�|n�&��!}�l%U�}۲[j�����f�d��	��}��c'�w0�"LI=�BG���"p�S��	n{�nq���Nn�cq����ӿA
ذE���W݋Am
�d� �a`׾�Hkrfn�'�v�����?rʌ�����q-�k?t�)'p��0����N�/�T�*}��R��t\�1h`;�Ж��~,��i�:Z���A��vü"�!+s��%Zn�C&Z���DF�F�U8T��Ϸ���/?�z���E�|l�	�ޗ�n�칰.�WQ�>ܷ��4$�Oy A�)HN�������}`�� �.�U�P]R�=��<�C�}�{3��^�Ρ�������*�r7�{Z�2�N_\�:�Pgx��s'E��ƴ,[ea�1����*��H4��l���i�	�<����0k�/`
|��}��vУT� �XJ)�En�=Xh(��0�O�Z�M$s9��K||�UYu����ڊ\*no=�p��][��"�ꓱ[�qR�H	�����.�y
L�����N�l.�ъ2�\4Ww�M�h~q8���P1.<�,C���e͑
����
����'^.R�Y�5���W�ԗ�"��[�!����G{M�:�D�t��#��Y(/VC�HP#N�-67��	M1��
}�G(Y3s�@��O(����B����4m�.ٻ2+b�����H�h)1)���$���.���kle�T���Gw?��|�[.��xsB��L����z)��z�Ǧ:\*%v���`F2�w��:G5�����}��bb�C��A�e@�}H��Au��P��Ȥ�H����_� ��x�
���!��r�3<Ҹ0�d����D��͒�G$�!~T�� �^�'��-���ln�3��*,C���8.ߏ�6�O�cXZH�c�؅Dg��tI:���@om�E�6�x,0��~U+~FE��i=\�Ҧ˼���q`�*��hv6�'�nJ��{z����.	��[���2T[��`L�"����S?�uF������[m���Z����p��ݓ���d��Q��z�L�i{����#��_�F,��u�G��(�o�*+���-mJ���ۣ5�����UP�l��"�M�$�eA`�}`����3C�3;�i~Ju��K���6�p]�p�^��s����ǠBQ!y�cB��L�4���U���˩��K@��&c::9�K�|37\ȉݕ[ߨ�;bXƄ���F��?Fw1)sa�V�	�&W���s������(Ba��D0=��D���BI�h�f4�
����"p��D��$��ְ�͸�S�oy1Gj��;�D�3S�����`�E'��ԟ��C6�c��s���@�3 �D��{
��I޺^�\^<�*�EpkTؕ��NǸ��G,�u3z�E.���DZ�D��!V2S`_���_��t���Lᜪ�r,<�+@K�0%��>e�����u��D��@##!��o�%AS�dE� �8�6���9Z��rVy �zD�zIw�&"HJ�7�ӣ>����Z;���Mxte�2[��
��p� �س�\���Ky5�2�V)s�IWRˉ��-S@	;�^k�~#��t��ӟ����g�����*�̮Z����3�Q���r�IPZ��l!��2��a�U&}���<�$Dy�m[�}<�K/l�{��_؁���.�ދz��<R,���c9,J@�;�Lay�+����N�+�)�b~���H.����|Eдם->��G-u�� R���"j�#�+ܺPY��U�O�-8�AT�5q~١1���((�kL���P��Y	'����Um3��>�O�@��/͋��%���U���X�q:�/��B�uvn��A�>�A�JT�sP�X�2�e�I�j�9��s]b2W<����d���	+��D$��A�Z��Yx2�S�[ǖtX���v5�KS��u'��� ����O�B��G��ҥL�����iN���va���vQ7v}y�L ;;��o�;�^��}���*��ڝ��T���q��D0V6���s��p�vb��Oo��X�|Z�7�8䙱*��`���mlx&��8b�n-�ߑD��ϝ�a��
*u��qUd�mj2�1�_˗Sh�,��� "	̕��eh~�@�3:��	bU��t׃�ƞ���������M������k�}��w^*z*?m�~9�}�"Idsn�c��~�Z�I�CM��U��!��$^�st[XQ�m�.��4�	ҩph�^����hr�>��22���̘w��aڷ�y_�d�Đxg,����EBE3�����K�R4{sK��WA��]��Z����J�@LQ��!U�FJ���d�Ӷ��r�%/j�y���I#;�y	T�.��M�~Y��s{Wrk��-$��/�ѣk��s��Ӟ��8�����н�3���k^�k��߼�>M�bg��(O2S�R��5'0�B%t�=�)���+�N�(���X��ڔ��hn#����Ng	Fj����bn�rpv�����t��ɾv��2/R�+<;Zg �����>�pȐI}�9������CCr���"�*���MI�#�f4�㾸06�����Ӧ��h׆`K`�?������0�K5|�O��Z���6U�s'���Y,0}�^��m� |V�[	XI��r*(7��g�Ko�b/�"����9�A��M�!�4c��%3�b����˴.��ۓ�e'�q^x��l�RxnP�h�����뤐�zV����C��(/�,��0]��e�0���,Pǟ:�@�zWxDګ�lt^�zl�����sH���8��T�qD�GiI��h�hbd���qׄ.S'���e�'a�{f��[~u!���\�����c� ��ڊQϛO�mM7ߙ��;�v|Š2��i�Tc�Է9�2���y��',���ŵ��xȆ�����u||�b�^�(�8yo�&k�s��+��$z���C4����n��\��b8� fw4q��pW�KZTs3��y�b\�ֲ�����j;d�L8���&��So��ɪ�=ZJi�gI�R���<K��u�����C�H��W�	��-O�Ѭ���E�x2\�*��q�_�3���$���y� ���k�D�mB�ڎЂ���λ$g�l�n%/����D+��y�rX���@xл��-rv�2u�6��U�� O�����a�N!T��}��O2em�˙���@y�z� ���uҫ��;�I?5�-w�z4n}�y�i�#u9���g�x�I10�=�)&��g�,�+��fe��쏄����U����ۘ�Q�\
{)S�ܣ�}T*�f�~j(�?��h�1�VIqE^]o�(�?Ե*�ߔ�W c�d����<'�/l��-��@Β��7�[ ��aT(\����^-dE�8fA�/��ɂ�?h���(%�'n8&э
�^G�1\��5�=�p	JL	����ԉD�K8ȅ\�JF2�KA��(1�_ݘ�{� &G[u��n��%�k�������Z�� X�ǴƆc*��bu��V0&' ���KU�8��w�A�3oΗ��K��B�:쁤+`�驈]O�R)��$ME;n��m��F/�H��n<?'���Չ�!ķ��	L�b$����7���:韮�KE�X�N���� �}���a¦�l���XF�ۈ�83D>΋^:4��G-��i��Q�K�-��#��7�Ꝩ�R���ې�a�+\�L��K�#����ǲ{����� lO(�����}d����m�D����S�+��ĉm"C�̯���z��0U���5/��W)��tU��	��>�x+Jc_��0���[��oO����m% �$>g�ሐ�wC���\@������k�{�-�M^Qƭs�Y�8��)v|+sd���hEx���t6pN*f��h�m�\�
׽e���j���������A�h\���$��D�uzgǳ�y1�hIC��D���\���~m)ZNp����f����llLm>�����g��`��\�^c-�/�ʓ��J�ܙָ�$����������J�� �����6E�^>{-�'^Ն�O.l��#��ti�胼v�u	T�oT�@{��?�q,�V�@��KE���|�q�����yi��R@7�9ްh�����~(��Nd:4�i`�\O�����*^�������|H��*�*3,��Ω;t�@}O�]���_��Tw���3ڪ��a�*���C�ϫ<�v�=.����Z&*5f�B��+�=DKK�(�#���2�J(�H]��D�d� *[�S�l��zݖ�o /�i��H�p�z���X����T2���#@�w�����O_�n`�:~3������0=�˸�h������qeS��b���~���ZP-�VIn� �Y�.a�d�4� �Y�ϫ�g}��e wU�K�οu������́�Y�<|�olv}T�6�]���m��A���(.Mh�݃O� &P��J7�H���A��6me���n4֮OV�uÐT�"�	�X�x���j+�s��h�R
f�����A���Jt�X+H��o7a��>����~�S`P����&1�V�9`���b\�@�q��wx�;�+(ܥ\��ڏ9�u������ĭk��;�q�������M헼�J��޽���|��."Ev����]@ۓ����Hk�2���b8��,�m���J40����l/�	�f�rB��L9(i�p��V�����4a���E�XZ�-t��O�*��7�=|��?����	��=5�se���V�u���ˎr��>BT�$��cB��<N[(^?C(�du`�8'kk�ts!��'hsÞQ�%d",��'�Ec9�\I�fJ��^�E��Id(�%���t7"�t�shx9���ŷ0_)B���؊7�����;��K�ƍ�������3Q#H�V��Ӎ�y��
q�9:dV�lt&����$[�*a(���O{A��k��V�9�j��v5�჉e��9IaJ�$gQ"aw"�97b��P�c��&7Dm�om�H�G���#��ijk;}9���z �ݠ"S<�����y�2�[%�e�Y �a��*������:剷[���V7؃�@p��!�m\�+I����0�>Q�e�z�^��=���>e���P�K�K"%�*���u�M�Xw�Vn��k�n�� z��ג,2Q��Q��CB�j�<��>��1I����uV�VJy��s��'���T	��N�|����r��峑�*�V�[��A;�j/�˥�Lz����_1CWV[��a��NE�#r�x�x�`�"�� ��u��]#>��o~/n����ո���_ÆT̰�� ��Lp��#�ٍ�����X(�l��y�ي���	/�4���#��!��{Z'j�3�RYF��l�3� �pEs�
��/�,f�I�z�����Ɠv�F��1�2B��8�}���E�ֺHӶ@0�*�syw�~N��i�*]����U��̏�IMak�,<^���հt �$��Z���Q/X�VX��f���	fђ���i�Lsb�A�ʿ�@c�\6N��^P+�����)�ncܞ����)d_r�ո�J�uc�}v�)�y�S��s@e�f�|��z���
j�Z�ZŮ����w����$rr����ډJ[B��Qg ���UD������7c�|�J`�;Ul��u�c\���~�J�N��H��3O3�R,o�j
�բW���'�������������H;Fp~�Cfܐ�}QA�~ �]�K�-^rJ��'�U1:�2�C�a�m�v�}*1XZ�rgD�B+���n"����'?ِTو�91��#qf6�q/u�`���~	T*��k����ӡ��vx�Ϳ�\�>j�u�����ab��!Me�0E�2�tA q�T�����?�V�2�iRj�Ͱz��V���a&�
��F9j-��M��.��H��ž��]������"�_I��w����ȅ���&�NB`��@3�9¬�)0|��BJ�e��Qr�?Y��6���n���޼*$�4MwD"D���}�w0���tP�0��fd��\A��.�%p~�ێ�!��j� ��L�Æ}b���R�;���>+D}��$��8ʱ��P���+Qf���n�h0UR�h�	�4�q?u����QG�:��K��r�X� դ�@!޲m�������'�#ʀJ�n���p�g>ڡ����ݢ.�����Ѫ�8d˃�;n�e$�d�X�M��� �Q�mqQ�Ք_�@s(�P.����_����|S���P%�9�Q�eY��\�6=dcʽ��{�h@%�\jm�|���k^n�J�Y�efbD�x;w���EP �Vx��U�q�Iho.�᫿i;B���Y�����ݶO��ºE��O#�w� ��r��3l!��c*���>Y��K}�yZ'8��HZ�E�,wƜsCB4�x�ja�o$b1�C��`�/Շ&�>�S���d��ӹ�|n`���ѐ���(��3���a�:o�#���Eb�&V ��o+݋�l���}�:Zm��[��$� ��ˊ�q8����k�.��U�bK��φ。[B�<�ڼM�Br~�^�&Q�]U�a7�tli��]���P���Ch`�	���A�1��L�F�\�bc����X��[�avp��:���-�w�.�a[�bc��!��	Ue�0�����1ή�mc��rk!qU:�zi���0�=�I���$����N�¾�X?��<=��N���E֩�4� �`;@�r�wCbE)~vY�+����I���i��ZдKD63�?�%x�.�&	��&��l��\���Ćڈ_ʆ�2_A���A��c����%!Hc�Cm\�˳^&%j�G��3�b�w�6�#�P#���Ѕm�;�,s]hƨ>�1��:|S����d�lDg}S�y�vq��)������v��'�����o�X����$.��Sd��k�=r��E@�%g(#Jъ�z�� ����q
��A�8joO!��u�IPFx���(_}ĩ(MX�\�wNcRj	�Iq3�����A4�f
�׆�ͫ��&��0�f����J���;n�J�w�{�vZ��ƴ�H�����_nـ��X��"g��=�D��w���ȅ)��%Y�ń�o'�3�t	�]W����*HrۯR�i\'�ϟ|69����=���f&��!����;�*�0�4A��~��zNq���퇒0����m��	(4�WC�p�>�̘@w�8���e�?�Eu� k`���X�m!A��éFzf�>�� �I?7�9_�9���^<�X#;6���٢�G4�3�4�0����g^�nз!	փ � �+�C~��=Z�����8��������#�-K�=�8jq���H��n���Sl��޿��O\������HVSR��W7�ز��-����-�rTO�K�
at��z�؉��ר�s�OI�$��W��?��J	�
��<��� c�_Q�=���i��vAW����,�=<��[���-�5��>"�<t�̓)IzN��7��t�}��
5-��<�	l`ڷ5�fh>�T�ڎ$����3[9���}L姽+y�iU��#G�O�*�mMw��臵&J�����H'�`�iixJ��́Qh��}�G��{�b��t'}r�((X�2�Ӏ���T�]�8�"6�o?�)���%�?p̿�BbH�䪟���a(F�/�J�%C��X[�`�J}�T�}��wl������4�q�0��:�5��'����9�D�#�cQcD�+�j�v� aw��n�r�Ģ�7�B��ҁ�<>�$J(�~-�r���ܼ�]q�E�i5�\�wp�sM�t١V�旀<8��1����Qxݛ�0wH����Ʃ���])U�T/���Es@� G4�>�㕍W*��@�2�	��(#r]aڑ�>�RW��Ւr�mW/G~Z�h���Ҥ���{�U4+�§R��Y
� ˀ���Af�_��Y֭f��Vn��E������&g$1��W�'@}���1��~~��Z�-��Ӧ�]_5�\�b�5B�;�k��|�K���=u�y/r�8���j 4���P����&>zfY�	�Yй��Z���Zr�g�S�1Μ�F�SVQ��9z�l�>��@���OӋ_�eG�NV��(�y#�����j���v��l�b�?)�b2�\�
E�.��&u�>y�@M߀����p������9�&9��^0���[��MOyw5@�vU�W����F���i *fS��ܷ�\��׻�G��d�l��"�L���~�f����MNa�z栊l-W�����bh62dz���8�1�ݳ?�Ld5��e�䃒��ap��o�ʵ�������d�9sHnV��Z��`K�����W�<���;�-�SzhG���I����$+IX��T3�)�Ɓ
 f�Β��X�;�}��l�k>*�c�1�m�"���h@��D|�J�l9��a��8:�lUg�i�<�<c�xɹ�+�j�_�v���pI.��i]�Ia0�m���yp)��D�/�~�����pM`��`���=#��U����/�K	y�M?4�W'��;�Hv�g��n��.s�v��鮓cRJ�a�\j��@�61d}j��tT0�@%�|�8�����1
b�+@5}���1�l6��k��Lx��d@Ήuн��k�*�s>~:��ܨ[��h5�m+R�\}4�&ʬP��,;a*��8�v��O��4�ƾ��>n j]��U�0����Je��cI��������U�=-Me%�ώ�nM	q��?�9ɏA�V4�n�'�2w�y�D���0txk0��z��K't͵߯e@n뎥?B.v�tO�!�>�hZ^��ȪZ
�;�M"�ŉ���|&?=�[���� |���v��Ȼ$�.r���5��A�љL�\n~t��L�(c=��c���&0��/j�0��N�IN�yw�v:�q��·�FA�9�ޝ߮`(�_����(�ؚ�u/��fa؍ƒ.J��&]�� �Μ��}b]])u��˨�5_�y���*�Y�����Q�e�ޢ�y9��hod���r7'F"��~d
�����84�}SQ�q򢯃��+��S����U> Ҏ���d5��K+�����;���W�׀q%Ƌ��x4p#Ƿ��(�W�Kw@#Bh�X�u� �*8�ue`�9������x*���kkx�OM����pk5������T)���n@��4L��^��CU��R.��{M�.����ъa�ߓ�0��;h*��X��egp�L��M��w�V7��������!�SY���T�y�/���Q��,��*+8�q=�,��<�����M�[i��foq�,�C8�Y�mL)x��z�91s_;h�����7��a�u�H��"�N�� ���&����=RY�᫜XA�=�3ݑ	.=���G��'<z�Z�$)Ś�ܙ��E��2���jܻ>u�e������Km�B�;L��i.tԖ����r�ܨ��Q��߹ujI��=�J)������ߖW&?-|�O�욋���|�Ro��gcր����b� 2@#�L��
�vmF�IN4Uޏ����}�k�1��,���@�߻�uw����b�B�l���X��Ѧ�b�>e��b�Q��������J�;�^��n��v]E�j���K ���C�����n��A@�$�Lx�hy[�LSiS��$ �{�򭽿��l�����ӻ�U��
�zm�o
۵��͈�u���8���`����>WaB3x�~�Q�����I�^Y��WF%��dF�(��Q�'h�ɤ�U�ީߤk��"
T�!7�<������ĳ�E��O��N'��U��Z�R�?^�r����M����>�y�O��b]�֨�r�!<��7��� "������R;����<�R���V��7&�������K8Q��uT��"l;��Lm��*��9Wޔ��9mV~�(
iЯ�D�f�7���}�|� |��Z�fFd��w��RN���`�w�,��������;�`	�(N�g��&�4ⱄ��,��(*�E�۩�S��'QV��Em��ST��J�\Z���2hchrV�U�C?¦=�U��JH_M���!���cCϚl�3�R[�K��8;�pt�?׃]��1����Oe��vf�]p��,l�f�W(s���3��c���z��|C�]�&��mBI��?�z�Z���vrq�}�?��~�'+�q��^Q���P+��%J�9Nr���;A$���{��О�՘�h>��VГ��a�!����QA�!2�O��4��w�VUL��O값n��D�M�5��6}�T�ye̗vuD`1�&u?��sq��-��z��n�C�4&ʞ9Ə�&�G��P��1#�}X8P9�����9���rf������(u�Ļ㯡*ϑX-c���P�2H�XLr�������LBg��e����W�̺=6nJ�Ɨ" �43>�"�Y@$��Á��U��r�Е�K���]d^E�D�s��8�%��)P�˴��͗h6�1���b\��FH�!�2Aʊ���k�� w�'�tĘX�����0i$����(5Q�l,�pU��_I�	�'����C���h̬;��aC�P��|�;I�UV�.��7	�C��5�Q	��7������y���,�D��a����Sҫ���|�2�&�˿[e!�t�Nj���6��[���P�K���O��]7�D�ù��$~v�7k�?P7.��2��Y�\��a �6�~�x�j��\�Q����h�P猰c����4ˠ)�����Ix��ve�~�xX��I3��ǎ�'D�0?����©C��e롙B�>ҥ��h�V�S�(�OE��^�[�5n8Z.p�2($����\�� �?5���J_E�R�;�����B�^ޔ��]n1�*Huꘂ��ْ�u��o}{��#����|7Ŷ{I��g4=S|�Ʋ�T�)J�T�
A͞��B�ݧآQ�|�G�.����,�b����4Mo�3�bOB�)�S�6>�˴�I:������H��=PYGmNf�۠��vu#��	�O�0��*������Z={3yB.X�H����Q�:���~�$:�,1F�0H��g_���䑕Ԝ� ������ҡ�L2�k��o\���1����j8��!�<V�'��^x�y2����%aG%[໇f�#��Oۙ�k�s��a�����D��Z��ȁ���K�$K�O���D�]i�.���_`����7�0�C�� �!���%-df!��Ə��N���U�	���#"�n��l�:�|v<�R硆���+=\�����۔w�vp3$<��2���V�ȫ��p\����a�R��\7v;i��)��F*����S%p���Ԏ�7�"76�Z�,����5`�׽fAC�VQ/ (�I0�^џ��绐vm\<�Wb'��bk��j�ǃ��J��.�p��l�_=tub�Q��wZuBx�d�7����}נ�z�_N�r�����^�y}]G-�A^�'WE�Q��qY�u\Xe��8\t���f�Cr��;a��2e&u6y� �>@T�U�#��b�t?���S�Yn��������XY����P�U�K��k3w��̿7c䃽��P(%����>ʓ�Q8����U_V�\�:NL+pl[u�H�O�e��͊��쥉���RI9K��r�u���¼���w{��S��V�뒽a�B���,�V(E��6�|�[�T�����1�%7PZx�4nMJ|D��6+�<V����dė�%^rs��7=֌�a%pQ�:ru�^�0k��C�K�Q�,�ț��6�K�ï�Ww�$y10H���$#�R��P�?9˔�U*廰�∗3ZbVg�yM�J�O[�UI�I�]Q<s͂ �!�zz�>quJ8_��
��̋�'����h����b��lݖ9�o�_�tW��n,�
h�ô�k��5����7����m��*���J.���ƩR����B.V��*���{�X����.FѰ�5��R��Mdİ��:����/!BE�>�\�Ԁ����Z���h]�(���L��v5�������t��}e|�49'�e��:�~ǔp���Ẫￚ�)�QFIs�c??}w��\�;��Ԋm�ܢq%�t��\Q� �-R"2
��;|ھ�&���{P��U֍'�iL�w���q6�b�s�����SX}>G�;�+ =}|�f�nB���Jg�c��&^%m~�Px��r���:�vFq4���lTA��"?�4��.ĂDO���:�.����")E�cm����Ȝ	m�Aye��w_y���dRZ��Yz�l�Kf4�I��O�5��s!g���l�,_����\�P�,�{�όM���M��uw\U[�;�@�/gZ�S�=�ZY=�fC%�ٞ�$7]�-�J���j�w�=I�$eѣ󍉕��/��Y��hWj��2W*[���`=��o�I�S�����o��*����^ ���(ND�l�0}�lĜ�v���|dd>������ VT6�7!�_ʊx�o��k���45q�o�[�2��L����.`�q��I�w\��l��eu�8`f�1K�ꁀȕT�=���ne-ә &HH�K��������H)��fxbvF�sHԥa�O龶&-����sc�ٹ+�����
���j7���sY�W���5)=�S��=n��´h�(�[�5Lj츈���}:c!�\�˦�dS�O�B�Y�VZ�:�{v3`IXs�ٌ�N{��l��!?}?O�f���f��U3,o�::�ޝ� ��W`���pD�$�$��wǸ�hs��˛ ��� K�a��-y��g�ᰦ���T�� efFHU�O{�:���fHB_M�z�A� ��b�lX�{oW�A(Ԋ��Uf�����C� +m�yy;��4�Dۿ�g�.z�^�w*�%�[sS�&��O笿� �l����Ƕɧ�T;��#b2����T>��"b�	(:�4�h����Բ���J��@����\��-8kaKdՠ�}�-�9�0���9uҀ�4�#�� [N�L��Y؟�s���q�������7��Z�b��2\]�)h��-J����_�T�9׷M�u����f�ƟS!�aZ�`T��TK&20c�@v�?��a�cB�;���e�#��u�H�����D���<�G3�����fCH��M�R5 ��+c��<lY�̞(������>Ѡƨ�MƘA��dR^A��cO!�X�W��Ev�X	|�b`6필ѣ��X�����_���=��UnW����6���]���E��}D]>��<R��L�dl��h�2�g�	~/M����2���d�m�#���0�d�O�:4�>��ю�T/�35�ֲ!	���b�C+�2��jz���"<�o:*��;���/P�"��g[
�r$/[լ.���_t�3-N�Φ���"D�&�@{�����l�|�v�Aj�,g�-aSǪn�n�3��Ox��Ձ�A�+4K��3��n]ư�l$?
L��i b��K����֦�,|�Z�7P"��f�l����i�A8������'�Ԁ� ��;@�ɔ��{��^��gh�69�@�6��YO[H��XG������6;�#�Q�m���ӯQ�l]��ǡ:f:�e ��GM3�W���Z[(vlN�;��:Z�#ݒ��܄��Z,j���*�.l&8�dڡ^��o���ګ󢉾pF=�s@������C��� �<{M.>?C����vf
n����.�.���\{�nC�y"�D����&�%���jM��`�K`d ����!0��H����������R�:M�ej}!f�/�Vä�G_ǻ�^���W�^��ts�P#���4M�vq�Hj��,z,������D�|7� ��)�m��%�o�G�G�Ȕ�]���u��྽���8%ʴv)����$kg
��6	�|�Xl��8��hk�Hs:vE��~��#�KE��ڽ�'Pǩ)rE�uR�N�m���!^�d�5	9�Ӛ}�K7'�L��p�θQ�����i�kd:�|P�D�(��$[Fp���$֝ӽ܏��t��1�+�T�jt}�;�#�ٟpx0�<�®&6���KL�<�>Ti�Pa����{���R%�>��ت�_�Ux��{QR M{����W�TK�&;͹ ���S,Sl�-����VI]Y�*)���=����ҫo�7�����H���?���A=)��x�"�?��)k��!)!�U���V��ے�
�>�5KL��m62��5	�^�.I+�
�к��x�v��iF�ε�T����ƭ��إ���]B�^�Md$�RI�l���C��$��`yyQhv�I���G08���ӻD��Z$�ȲK+�)��mSX\�_��� %rԪV��� ���i�L���Q���j���H�Q�Z"\�(Ej��9���>��N�����#;������x��h�J�;d�R�$�:�R�����1�����r�a��⌴.Uط(n����	���A��@�^�k�JF��8A�Pzޔ#��'n��`Ɋ�����f����t1�T�T�'t�s^©	O�" ;b�CJ���$-���sQs"Ӗ� �>Mh��]�jW������;Ps�r/B��m<i��:����FR��o����
���S��&M�Q˰��8Y�Ϋj;d�M����.��-�t~xơ�kP-˺�4���V�?O�����`7ָ�3�Oa�*s'\�Ӟu���rQw҇�>�"�A
��`f�P��,���*� 2�lECbJ�	E@?�l�a�mL`o=������ڡ��i���a�C�L���\���BP5@]d�i�B����Qj�	��3?
t�}P���6���@�E#�~5ygZ��Ȅ8��z;����7-��b�'��z�����������e��x��S����ȗcg�cw%	����&�G�5��N̨�`ޏ�.��.��������RX2�7����6G"�]gŬc%V��*W�ѳ��SVu��}K�E9R��OЪT��-.Ó}��Ne5��ë�4VˠQ�gJ�|���vXM��9�E����e�D�-]�����'�%v-�l���Mvdp�tM�b�_�=�@zN�hFu W��d�nv����`�����V?�n�L�1ߨ����ʰ�ͮ.��"MUh/	��������j��B�n���Y����:Y�d���� �ts=ﯫ�$[�`4��c�g,f�[�r:/�C�b��7x|>_OH�h`e�5!���XA{aɳTZ "p-���"i�HwnH��[Gb.Q�@�A�]�ם���S�{D���~�M�|�utk��-*g��h�%�Ny.Hɰ(9���9/�^'+-J��䵗fVB>S�ۣ��Yg�ɼ���ؔ����<Wpi(�4<P\�y�}H�k�
�T�=d��]*��J�+�E	���W��{�!:�O�ی�'�& Ŗ���`�ߴ��Q����o��;�7��ųL1'+��:��=�����rf��V���(����;bi#(��'M�r&�/M5�8X;�z�|���Ђ����:�ϸ'+̭-p�Qɼ#�t��$��*�����O�eP�4�x���g&�-�*K�4R��:��Z>�$�p�r�ށ��5ה��7~���[�x K^߬Q*(��H%^�cl�_v[m��G^0����1}�Āz�f�4��n�c�K&��U`�����U�1�����
R&-ET�[��O2�4�k��mUԓ'��=�YH�^8�,O�T�Ȟ)l ��\Sav���O4�{�{S�  �l�}e`@��Ƹ�^U?�0,�<f/��}�&�{�8�$������G+��9����,�k��Wp7�,��8� ����0�b�~�rk�߯m��Y3���c�o�+_��
�{�_ ��y��~�b�z�H�I���׸;�-�.V1�7�q�@�����٤&k|3}mUrp`�y���3Ӓw��ALzˠ/�z�
\� �4a��ʵ+ �蒯�ج�rY4j���|����C�Te?V�e&��J�F�A�&��t�]��b��eԹ��!fhJD�;k��¨�惤C �xmm�@�V ڠ�iA�ń=�.�N����%���cw�E��"���oj:>� �uD� �\� �#&.�f���ns��d����|%��Z	湲��I���H�L��+�����TKu�/y�H���ji���VC�'sYN��BQ�&L�����F�!>RWe�J���ֈοt:ͤ?�W��J���;�۽�x�5Mĵ��o��[ ��@-�܀�Q8у�����_�D���� ��;�#�LM�̊ߦ�Z&�G3�˄�E<�m���z���A�v�G�+�~�G��ͩP����#���\�j\�*$�=Y��`�#�B�d*�O���!!����r�
5�KUB�2�<s�=�0a� �,���/�ޗknI�(��6������pS�5�@�~����Հ�,ȂF��P�L�OCh�?p@���p'
,4��U�c8V�z���d��1�\��-�����j��}�R��Hܶ���$�J�$���8�E�0��Y�{���bߢU����ő��%ȸL��M !��Z�'�����ynƨ�A�]W�o���2�7�]$�m�R��)8lZ�`^FPjv\L��9D���=�����	�v5�T�^�'��,�皈YG����k�H�%���*_�����@D���*��¬�^u=�Pt�g�JN�&�����)�_e'�ǥ�4&w_�L@��m�� ���Z�<��Mz&�����o<4f���r�;(^�����d��-�[
j���<���9��C9��U��-�)�Jy���@�Q=t.�����̸��g'[�G<~��gI�����i22�+**�1e�)�j������9K� Ւ�c�a��L��f���ǂ�%x��Έ��~b9z��Y1�Fc(�<���>T�j%��^AMŴ�w�@���V�_;���'�f;�{��VLu�� W��!����h\���u�HB>�\��'��$�B�^�"�4/��:���������1�lv��I�<������Q��8���Ŵ/�3v��_��%�?U/�hI��a^Z�$R+��&�8��J��QNz���w�5`�ҥ�w�<�{&򁎙-����}�>�|S&>P@:ң!���F�d�����`-ì�X�2�1�QU��G����Aȿ�^O�L�X5��}m��Qg����R�h׽l.���S�h����ٻ�e�r�T��C��i�7:R�_B��gw�$N��U�Zj������+�K�����I%��L�wG�;�F\�.�/�O��kI�͸}��6He ��9�ɦu?_� ��-�o���O�5�N��\���a�U��ŠՁ�z)ϡ"&�U�~ٚ>"����L�j&��'%cQS1�n
$2�ðbZ�:f%��'�(*�=B�ܹ�[X��ПUGb��/��F�3X$�8~�V�p{iu,��wZ�<I �+�-\���~Y⯊����0�ڑ�ܜX��B�E0*:=�2%��W�+}i9���v�LAB�(�M�d����3��k\�g�����
:�KiH�2�Y.�B7ט�qH~���Ҷt���%�%	�%��3����H$N��^D1:|T��wܜk�y���U����]RϚ�en�G=LmV�߃�O�vv����:��4c�F3�M���ݛg�Jf �7�5�@|zXM�-���hu�h����K�p���9�����a`!̇k���i�q��9�C��OZ�᠛��*/6x��3����i����{�u)�8
��F�r�}Wf���M��{Nyyv���-���H����V�F���r�T���*��%{X�zR���z"m�/��%�5E����v��^:���,@7�쯺]��{Ϻ7��J�ƀ��,N���@����/ƚ?.�u���FK��Z����	iGM
.w[�➼�TRZ&�<�������볃��v�~y��g��%s7G�KG��z=��D8�����}�$5�2,i]�$}\<��>��O �!N��*��=�ý��i3�;��CE&�eD(J�m�u
}5.��o�� ?�+�V}������������LKY���ԙ#���չ�2Y;�:NV�bz}d�-c�;�5�_e�j�M�kB3�m�FvU'wg�|��hR[�_hZ#2j���c�D!���`мq����U�o��I���t�	�r��O�#���,V��j�z���Zk{�̍�g����������I��u&En���D3t�g'�������1������2{/s������9�[�~o8U�q'G�P̀9Sҷmr7���7`�T˚w_^Ο�U3Jo����O�9C-���Y�\pi��Z��NPA0�=����MoE�7E:a[�R�����d�ri���ɥ?r���R�HN,.Vؔ�ɜ�w -\���|����S�ܕT$�,�T$��];��A�f8�-ia�U�7"� �e���\��@>�/0�����YXO�u.�y��=Qu�N�,�|QyEmw�(�&$�!�4�N��u�TSڲ�
��cMa4����I���"��L9'�M��(�+���C'�����ևu��:�%���<Xi��萋�U�]�_��cN���%h�>Z�r���Ϙ�J��'M�u7L�V��h��o��N֘��`@􄖽��I�T1!�N����w�����=)-�w�Oj�84�)9���Y>���/U�F�/a��$�^��b�Rῡ�ռ��$Q���L�1�h�M��!�f��i�]Y׼,%"��B�� ;l{��'��A�ŗ<+�dt�Ok� �r�]a��J��#r�ߙ��c]��2�0>$i �ܷMa5쫉��d���q��R�W3x��fo�.	��)��UЕ�^�" ��RRs"�aޱ���߲����X�]���w
|,��l���P��UU�P��o�-!M��p�S�57�U�owR+�E��Lwr�f���w8�O
� � ��=����"Ue"�#���?�޲�S#2����|�̝�+���h���=cDF�4�(�*t�����6l5-l"��I�R��<��]���쪙h�GMs�'�M�B�yh��r ��L�k}i	����o��ŔR��/>=-�=0��ia9n��/'����=	��پ�)��>��|���zk��TN�h��?"9Xѝx�ʩ�0f�5�y �Z�H�Y��}-����Q�D, ��(T���J�ǎ�/�����'�����#<�����"�x� �,+�������c� �s�1��[������ޛ��'��SpFX��F T$���ZN���t��w	�(K���9Hu��'���Ⱦ��և����Iu�D*�͒��3�g����`|�-?�-asÈ�-�,`�m;�˚Fq����LJ��yҬF��sRy ��TP�#.BW2��>(��6x�ԏM����`����������l��&&�{�7	�i�����cX|	����%���j��:�.G	=��O�q�(BIa�z�2�CR�hT�J�����	
w	4����\����Jp�[���i��6�$wu·��: :u��6O��{�3Q ]Em�]ܹc,�	�?�#�	^����DG$+�,sӧ$��@�f���`����Z�s�(`�uv�8:�ɭ�%g�O1��f63�g+�>���W#ioQ( �]i.:2� d���:?c09�>NO�I�\&z#�\��m�?\���X!{�1+dj�!=՘ h��$̔ �
�R緧$��5)�6�61��z;�4���փX��QzBL�y�,v�ޯm��w�ٹ� O+Q�?�f9?����1q���fn&�gП��:U@0�~�c?��홡�N��#���܊�ꜳ	
T��ln.kSB�M�Ux���<���q���%��8�RJ���J�r�tT���h���o蜛��ѱ�.��;E �쵦b�Z��� �ř�� ���LR*�m� {_�oŇ���>h�I���m8(�@8o���A�4!a�F�.]�i{� �JϪ����W��8M<UQ^�#�k����K58��ۏM5/��`�797�D���������;�^����ͱ��Ϝu'ͬ��z�k��2�})�����S0f@j5<٠L4���o�'��� ��Ic��=���~R�LxP�9K갂��D����ջ���A�� 9}��@9�^���Ikiy���4��gC㒲W�S
�滳-:Y�DeA��u���^��V���r����/��
����O��v
s��7�k��![��h� ��K��=tqMƏ>�:��g8������N�a�ې�(h��VR�{��zY���T�Rއ��e���7hu�2<wJ��}�?aD�����*'���Hj�%c�F��&9^��R�&�O�cꒋg��,ؚz&Ur��W����K.f�?��j7�c��s%� #�P+�w�4,�
Uk��2�Q�=xܿ��հ�h��e�wT�d���=.Uat�g�<�W Ӎ�c�d�]�~�`��8��(S�U�
��a�U��B�`~��5u4��C��IAAM����a
���l���*:!E�M�D���_�����/͊�
�ǃ�>c��!g�]�D[pKg���Z�� g7*�C�(�7-Z����w�߹�&ߨH�B$�]	%�-��&�������sW�
���ҮYD��V?7��N����C1�oP^\��gVF��U3����0�*(E%�����{1�TPƷ�����^�Y��
y���R�1���dH���1(���]0�����8���H���F�����^�"G��!�� ��o�ԛ�.J���d���gt��ں&D{(»���,P��oC�]:{�uu� �V�H想g���u����@�D�W:����Q	�c(�%���f���O�]��ES��nU-`^�!p}��/Vġ���L*�����,��7����)BuV�mO�%Z��^�W�z��)�#�#����n�[�D��� }�ą��)�)��H��.����R��R��-��9���.�xS^V�@@�66�V�9=dD/?.бY����]����vAJJI/�(>���ЙT�M�d�Q���tu�%��X���	Ĺ/���c\UW��/�
S��C���㍔������x��h���0a��V��<R��P��mG��B�ڳG��\�:n�����`��Cm�^��nJ/]�6���b+yqH�RaQ��:�����X&��K[Q*�A0�F�|���$����Ӊ���U;�A���4& �$��Ld���n�Ǘ�I�"!3�x�1���j���kGp 8yH]g�]�w_�+0�N��6E<�)yc��<���&Rzg��wVu����E|%g��حf�!k!<�]f!VR~�P�⮘Z����a�¶��-���)ϊ�mQ����g�d�~N{����=�mʁ�$��:��Vvr"�D�����Ѓ�M	OA���x}�\��[�=#�z�R�9&��+�x�*�
=����ª^���D9����v{.k����PFspM]�_O%�r6��}��/�F����Ƀ(t�O��A�����D^qʰ{Fu31(����-��Ҩ��QP�:��A�Vk�[a��Z>� $��?�7��l\PФ��J��M����ٝ;2���Yr� 򡛞<��� x�{\����Vzb���ĿA�Ʌ�V��;E�4&�����di�J+���Ĺ�g;<���h80� ^�r�o������&NX+Z=z�B9M�CC7�; T���fg���	վB7��,?�Ow�"H�W�7��X�m�۲��D/��VƘ�ぉÈh 3��A�=e�4nx��R�ZGU���a��R@��P١[&�hx�۞݅Ѥ?�0H�`��Ϩ/�M���]��W��h��S�nt�(Ƙ����W�I��5m�Svcϛ-�����H[��UV�OD��Ee�|�	(A
N�SE����Ͻ�l���S遑8d!r�͈Bu#�e��2J��r1Eh�D��x�_Y�%����Ռ�&��$��L.$h`O/��=�ϭ{KmD;�1�%���sP�����s���\�c�� o��	6ն{�J`��(��||�p�4ϬT��>��_�Ȼ��2�s�ϊ��:z,��2�M����2�t�(�&���k,d<F��arҲK���0�Vɜ9��ʹt�-V.2���qi;A�I�g��	ڬ�����;�՝�\_������1*�l=����";����=x���	��$Tn�	�T��z��%$�٨��h�Ǽ���w-}P�? q*l���6�Tc�m�N=ب�a��Mw��*|�c�|3j��O�d��Q�H8�i:�3�Ms�.���T����a���0��8��Λ`��k�o�û��#�_5H�<Կ`�$�;�p�(��Z�tڂ�jԲ��%�o����ñ���)i�8���Rz���3�t�"��vX�<�%�Z,;�C_�B�N�|"m���G�����Ğ߸^�K�@SW��l�$��<;^E��8�m��^���*ND���هo�eJ	$���;Ѱ��5A�9�
�R�d�\��<�gq�y �@�n��[����M�GĖ�?>-����kƱ��!�o�e)�T�'�xb��
uB�<����I�h8;a��ñl���!��5��A�H2�M���T)h̜������+>�"�Va��/�Z���-zڪH`�ؔ��[���e��[���j9��l�1�y��
����<��������h�D��k������ml�<}��Ĳ�'ზ *Y`9U����@�ܥz1�s�Y��ǰ�Gf�@FY�p)nQc6&�mSC���M���
�E]R�G�#�$Ac���>�ҁ�E1$���cvùc ,>���c�=fSZX$+D�`���`������7 �t�Z��p�����F��oɚ��C�pܺ��S�Cp8�|��4_R�U�;R�\nC�B�/i �à��㣧&ig���,�t�bn������]Fg��m�}�\��?�Lh:��}n~���RlJd��?�M�d_-7-pZ�R��#�v͈�V-���W;2NP;o��j���A�iԫ�b�pGQ&��m���a�n�(jQ}d|
�H�JG���4�ve�<j��3QA��Weh�|��#�{a�W�;�Z@����s��<A2:e2��+��/�p��O�5���c6� ���?� ܦ��������i�O�\y�H��*?Nʆ1=)�	��W6I6���E3��ؒ2��V�66oa�8�Ա�E��2(�%�8R{�	u�����}�e���{]�:C�;F��uW�G�V?=�L�X	D@o�����|��Й�RÌ��;�¶���bI,%ɘƘ��IKX��h�:X��g����>�ɜi�gv���]����T�ј��ǐd�0��$�T�.���~-utdc�z}���y�
��9a����x��A�Bq�=Q�%:�Ce\�5���A���B-��ħa	�l<gY=��a��"N&���`d��l��7R노V7^P���ȵ������`�0��gD�����3Q�����a�Ai���jwq�m�'����Ḛޜ	���$����K�u5%�^�1�����N���έ��I�;˞v�Z�aݍx~����Tp��Kb��g�K��� �Gd�f�� >�c�/�T�(��<v�Nw�?�w �H!g{�����M|P��H:b�>�Z<��n�� ���M�[��;х����oH���E��i��:��qJ63����|%^����ɠD4	KnE���9��0Y��}h�9���&\�Ĵ�h�����X=%$#'H�E��$D�J���e��Р����SzY�%�<���/'�u�-����b²��s��\�j$�, "Ƞg]f� �-��z�⽮MB$0�H����j*���m�fS�N��A�y�0�dU^;.�A#f����p#�O��߱�9����O��%Hb�1}�RWH�c�}�v>ȱK�y^T�td�B�&Z��F�JP�9�隉���&4�(j�8��/Y�iܢq?�t�n"�k�!#
�Z��,�&0�q긎�G����UFic��ʓ�BE|>^��坲�D�f���Yn%nQ�O���zdh���h�I�s�c���3/�ʠYX�KQ�Fu|�)������B0Q�d��Ef�у�2zMB+JLt@Dj��k��8궰�F�T��՜ʜD7�|����cN8~���6�S�<��v�7��F� M���|Ն�j4q9Ki����ly��4E�c1��M::[�������#�3����zJ�Tqbj+:�8����P��>�� e�1o4�D���3H1\6�,�z�`Z+�ADÛ�� �+�S�w#��>N��.�4�!��� ��Q`߁�6u��,*�����-,��GD�I �sZ��	}B]f��z�"	F\�����M5c_&�?�i�S���V)��+�?�@�* N;5��`2�ԧ�%S)�L�WԐ�1��ܛ���	�$�1��Dp���%
�|;�����4j�{�h��/�_t�b�ɋR>x!����`����??��	nGE�l��pِJ�	]6i!>�f�Ds���-���ߢh�����Zx�Ζi����(�-�Kd�v��^q`" (��\�aה�1?,��9|&�%���S{[�d臚1)U@�6h	T�ANf�E�E��P�X2u����y2�+!�����#��(o�����U	������?X����I��)zQO�{<C~�N1P�%�!�.�|7���.(sv�4�����q�q,Ù��a΍����u�	���{5)?�t����{��?��H�	��uHPu�ۖA��m���',���M���т�^w@ȗR��wD��	�c��R�_ϲ*�s�j��	���J�J@�i:�L�P�/>)�\r��ͺ�?<&����nH�D���iex<���]�P=�"�AVS��\G��S�:�ȕ}��Q'��ɪٍ�~E�&�N���2lV��2z`��+z�hT�r�e6ÅՎ��x|:�(T)ۼs�Ů\��Z�-Ln�R�E�<�{q0|���yBK<Fy�{���(%��m���rU�ls+���'���s�֛��.������	���sU�����֔��T��`�Й��1{*��s�5=���.��v\�Y�:e�F��M��/�$_{�]ܺ?��Δq�Bs�����M�܊_p���ia���	����B���"��+k��<*89B���p�b߻<�o38@b!Š��L�ɘ7G<jg��N~�4�C���3-�^�隻�b��n�ư�I(iZ�u�l^�p� u's�wO����U���c ��i-.Z �Э( U�X�⩸��8T�nՍ�n�k+��s��FЋ��n4*|��[��GoelΓGH�l���Mo3vD�QC�m/��M���2oJ#@G�8��J)� �q�9�ƌ_��n��ր�0a^'�v0�q=	:W��w���+Б��V&��9��m�`������ܸ���t��υ�#���EW,G��3��}��heS y�}�V�I�*C#�h�<�t}=�Ɖϗ"I䉺�j?���M�:	�6�����)E�+cP�8��������>��s�R��S[����E9w�o1YI>���Z-���UT��AA�Q{�=S��M`Q�c�%_-l�K(/���w�ZhX_L
`ӈ�/P�f���c�q�-� �2lg=/�������Ё}<g���;L:hȹ�� �R_Yz��|o�:�k
+z�S���ׂ�w�a[�ж���WqM�a�mчh��W�9_Tʎ��G�6g	+"B�6��4kR�J)ʉ$n4��d��`= ���:��$����Z�袓JF�^S~.u$�pR�+Ҋ�Xʠ`�ItDO�|��vxZ��gq+����O����E9�;�p�Bj���tR�.h@�Y�p�m&��	d.��<DC�BA�}b\���c��T��Ȁ��7r5I{�8iY	}�Y�~��^�Y�{�_m/�q�|υ3�|`��c���%.��;��]��;b�~j�mc�1�)� _l���ϑ3]�	��!����d��: �Hլ��LZ��Ȅm��]Б������x�W�!-]����M|d��Ky�s4^���@+щh�i�H��z�w��>��{����{b���\�!_V�h�%�P�_cԜpL�t���a��Ď�������z� ,�!v:��.�U�D"+��2�(�UY�|��m=��,�ژZ�il<��]�z����>z�c[��õA�0�:��0+�.�qwy������bߍ�'�M�\
�n�i�6Iَ������<J �QR&bڳF�z<�A�[��^��G1��D�e�G�qT2�Y��}�8�C�ymG�� �Wp�\~���;��:��Kp�3���`��Ac�#���5�y"Q{(�j����b�V���[Mń�K�^��R���~L����xمr���Ý*�?�&'n����nP�]�7
e�Ɗ�O��� 
�G@��q�����m�Rm��l�&�ȣ�7�0<5���3���1�XuD0Ϗ��2
�R�j߁���"���x�Q3�3���d��h%g&��ls�A�V�*�<"���
��0t���-��M�FK:��z���`e���FɶC:ju0�a�E�}���ݷ<���m���j�{%I�Y7��%�����<r)w�Y�A����Q'�<�$IVf�EH���g�?焕�z��3���ɐ!ypsۨ��a�����0#�a�i��ae���H�<��uO�g!��^`G�ΊBn��$�q)s��:+���M�;���������]�z|T���1�	�Rue�VW����E*�M�CcpY�.������u�u+}�(��Q�<�e��a����/�̢�ȿ�H���7P9�L��bf�˥
bd��F���'U�BFrB�=�Ё�{Q<!;on#B�x�2��%g�aB����-���<�: FZ��0V��3����} W]7������=��>��US�������՗��&��Ѹ�7� �~�@e�m��F�rB���5����5SX�*+v�<Hu�d��֐��'0�,-���ԧ��0���'Lc�)r�x�XF�*��l��f+��j.ou�g,N�Z<C��d�NF�,O�i�	�n�+�e{X����>&���ߓ��ǫ<�Ew�q��g�;4��ocJ��z�G�Lȏ:;���2�0;�Lֱ�~���?(�E'��_	�Q.�;��?zH�~�_�R��uu�c0��S���'4G��?��\E�.��f=c�-����1�8��֚��"��v��"u����V�T8s_��P�������i�-9p���p�&�ԕ 6�~��&���B�+���o�
e6a�a�
ɆZ��KD��v+�[w���!qg*ٻB..C��[p�z�n�c�TvኃZ�3�Ob��|��RC��5��J2Z�ݰ�<��lΈ�Y�����A���|)~����5�����Ď�!aB�X��FD��0������7c�����s5��##�9�lJ
��-rK�K�(���y����k�-j?=?)?� �m��_r` �%�a��]�lm�H�[�6{�.�S����*�yO1^?��BY+D��L�����D�mv�3��H��^g��d��E�]̜~^R��9���m?�э��64 .��B���L��,��J@	`e?��z�y���������V
YPL����JE��F�#[6Nb��-0���d��>�iZEoێ�D�E#Z�L����-S�[j�6��������}���M���lnCC�P[�<���O����O{�R֭�=���	{��"MM_�����%�Ӵ��;bc+Fdᢁ��b"���V��;=T�l��Fl�N9�َ�������Y&GO��#�����HZ�ɾ��:�z�<���?~��D_x�`B���m×D���ze�M���S�*	 �g
l�y���`��x���N�$}���w��Tfߟ��3T2��b1EQ�&ވ��G+���b𪸋�xj�!�	la�bR���&rp���þ@��)��'�V?���@��Dx6T�XL���.��9ɔ(�/4�������ҋ��_WU��r�R>�k�!Z��?�n(E�~6���F�i_�� �z�����އ��:^l���ㇻұ�� q@χ�&�b�%��M�R�16t�$��$X�`�ϻ�Pg�1�\��~ ₗ(n;X3A@�����R5@h1 K���AD�$gX>�������"�U���t��ϡR{_}%���+ڒ�ë%�(��M��	�.��ɴˊL=��AdL�d²-P#t�d�_BO�[�<^�a���e|�r����,|h��6�5�,B�H��ڦ�w�B���}_��Sjc��8�c<���7Kڧ���|.P>N&T�.9� w���5"���(��;�b�=�������*ě��Q��vn����m�֘�G�t
VK�	��� ����]BY%A�7oV�mpE����A�,CZ�>���p1���~+tg|�$5I,�k,�w<|9�+�XZ��E�/���'Ws�=�dlf�+&����
���=�~�!��x�V��8���ԕ��%�.t6�mU)ynh�����P}��ؒ�p.������5��"�"�?�eIȷ�v9�Xv�0m��a�#�e��[�����������=�YHly�T闎O���i�0*��Q���ΓU�DfF0� Δ<x��:1b�߀֭�	F�Ү�(�u�z�?��JZsqm�XjO��K@;�Z� ^b	ɻ�͞�{��S\ߨc:چP�Ru٥�y��@� ��W���J�<9�LO����$�|r�v���hE������k~���܌�;�7�q��4��=1�?�a�L�}^{ʼF��׭w�Wy�1�.:, GL�,����HL�Y�y-�b �~��{/w�;[���KV��<A?����e�z���	�0�X��!�f�.��(���v=~�{3��AiX��8�e("m��_�?a��Z,)����#�}AغNu�Z�7�^`
��v.iHJ���u�,}{��U����ص���V
���E+�"
.�>q'����r��o�&�$po�34�Ѭ���Nv
%��5��F�b�P{��o\���S�������l*"Vǰ�7X����G<i>�I��F� �d�nd|�x�����dD� ����.7ϼ��e���_;̥4@K,C<��2Y5�exf*�=N�(!���!�{�@6����~�u���(e$6�Wx��R�9q;z�1���v`�E�����%Z@v�ağ�Y��w>8�|�Z���D{�|�n�|W&�J�M�ƤQ�e��U���$�A������qѸR<e�0�G�,��W/���:b�7��/�[ AS>3]w�����b�p��-S�/fO��8I�X;�/��M�+���X�qZ-	Y���=���g�ώh?RBR�}$uԁ}�=���K�t�ׄ�|�}T�zլeq��^����3	n����;�Ᵽ�N�}��	V���"}�!���J�BX�`J����8�C�P�2�5|$ؐ�f��S���huY�>�`���.�Hf�$�_� x`���\I�UpU�2���L��I�5u�s/Aa�H�P�B,��T!A�أRe��Z�6����D8&�ڝ5[�}���8q�P���F#�p� ��v�+"H���&�r.V�; E*f�����8`t�s�6� W�O��R�V�bʔw������ˑg���ٻςM����?�@yHһ������c�c��mV ųC���4����+�ZyfW<N9��I-!�C���E`l�~i7�.�,�~<�h��W�Dn�i�Բ=ͻ�i-�i����A]��执	�c��B�s���Ԩ�Z�����5W��𵌍�cIh5�
�RU��5�3y�z$,��\q�eúy�-" �-�� 
af*\g�X5_K�����0��� ���k+,Whj$�x��5CA���C-��Cw��Q~5�Xζ�2y[ZF¯P]v�^*-��z
�6�'G�aX��?�Mޥ �iR��0�;p�]�P4~ۦ�P�ؿOh���3"�<a*����q��Y��k{U���(��� �GIM���Ѣ��e�GQDLͲ�&� �f����Q���຦���0���ٵ������77�V��J?}a��y������c��V�:ގ�����g�c��.��wy�n�(����}:a���De,�~��Ǧ����v�_~�n�/L�t����!�=姚�����ڢY�f�s��u �.~�������xL�?�?��9nhr�>���]=k�ݧ��Ps�,���j��\��~V��I����-�_9�)޵�ō����5�a�ҫAW"�M�q|���T�w���:r)��S%(�T�c�[��F��h��k��c��VyƝ���ȗx�e:vw���#<�)	(t���g����(���V�o�W�5�R��V��b�]2286a�7��ё��2��[=��'�Z?��\�a�HDP!V���3���$�I_\ ���F�o)������0��CxnҰ�'m�s��F};;�L�`�C�s��b�8�˴�=�Q����30<E�����Z����Ɉ� Qc��/��=$ŉ�E�Ă�ʟ���Б4���e�88�����D���j��R���u�2�u�j?���R���g=�[�:]�KkŉG��S�V�r�;*��jJ�n	��:�3�X��~�19�Y	�#��3?'�2��c����6���Zm��qn�(�� `����RF�Aq�x۷f���L���O�N��p¡G���\�:��p��V�������j�X���pa����-`i8f�6�O\�%�ml@�x��i�lbW�0#����Tm�Kk�s5�k�:�r�	b�H�Mo@f��$sx$Yu˥L�����~�X*:�>����J2@�Юr����7�v�NK\��M*�ޞ)�D7���LT*���'B�}�3h~��D{ߧpe[gih(�w!�fC%�_S���Z��N�I�v�m��	U��P~
C��<�F��67.6d73<����JͥVT��V�����
~e��/�-����lL���Z��&��+�H߃�
�B2c��-�H
y���vFW��n���3�$�i����Z�����*��wA�˜{(�|�m�8]D��o�Ѳ�s�����J
��d�0�R��3d�t�bDWᩏ�ێ#�2�E��gv4g���{���D�!HpnF��Ď:=Լ��ߵ�B��5I,!~6�ʁ�s"�����L�蛔��;�4�p�Ȓa�q�׶`��}Cd՟��!R�:�7��*[�Aa��߆���,�Q�/�r&~�܄�zA�T+��2��%��P��|��c���ziO�2EZu�?=#x8O�[R����_��U�	�LkBa���~s�z0;��Ř��.F^u(���rpF1���I*`Vx0�?�h	�~�Fq�lQ}���lr���\�����H,&��?�FT��c[�Й���m�M�g&=��X�`�sXF.�t�z(�=��/䷶��0� xRc��N�<q�����Ag �a	 ET0FA^�Xs	�[��G�]y��"���s�|s�M��S�l1���X�s����ݦ�As5n2`�Ϥbwz�@.̎j
S��c���FG�q&#�:D��ݱ^������l�'2��x�XO��~����1~��
z�lw�v��y�U>7�m��M�޵�:"�Į�n�Ã�yC�:��N������>��c7q����G��m�UY�!"��0o�����]��[��Թ���h�[#��e9�XK{����{O����(���'U�y����Y_w��Uyⶕ(vi�gf�!`�]�.I6�
�Ԝ�1S(��c̆C��Tћ*:9����=h.8�w3ǝ��5x�+{��;���hs�v��I<��-J���
3��1��q�Yh$�]�g��wx�\I�A�9��l��ڄ��R0Xc%���P@�3&��0]��|��>�[���W�I%�m��OB;��ݽ�����d_z���,J��<�8��Z���H(PwT�����V�(�`4�z�2�	�3*�VL�>�f��U��vS!�L��5l���r)�z���E��.J5r�����(�gfUo�B�0����9���Rc�rX��.��	C�sQ4�ʘ�d��=Zc�)�N�L9�T����
�|(˭8b\�z# ���|^��iI����1�χ�����x6����.����/���ܸ�o!'��)^I���/&^��T�Nd'��~�>xUg05���[�Kg�~�M0�և��/?9�$9�_K��׀8;s��@�����؊�ղ� �S�`��G�M�H,����4��}�DEe��3'Rfn��K�7���)��'J����mC��Ѭ��%���=�c�?\uv$���Cdܖj��zE�H���U�n�p�o�Þ=�%Z���oCA��<����TX�.��1W�Ur+{$0Ԗ�!?r���jM���gK�y��^�_���� ��o�s]�"��0��z8��^DK.�W�'<����9��@�iJPGﲔ�e��츊����L?�LՋ�c�z�	XJi@g�I&�u3�2�^9��D'��%�+#AoRb���e�L��P7��D�~����mau�����;��{N��!��0���1sm��"L$v~xN��Wl1hq����t���9�0�0A��9�4��^�M���SоJ�h���5cir�T�A�}�	8hB�8J-��{��N��L���s��?&�����zlQ�@��%���X+Fm�A�
S:�@<J�D�9�uo�Z�h� w�x���C�NΆ�*_������kfF��#_=����V��y�"�B� ���x7C-o4V�7�{NV�C��TwO	LS �	�yF��r(��Ը�=lW�t0�p�a��W):[4��-q���M�n-��-���%�������bx�n-_��������~���Uq~�s�<.���?����8v{��H+���ܬ�⌬��|[��#����J�Ô�;�C�o�JP�JZ�f��5�[�1�:���T1c@,����S��Qd
���_QQ�����ߑ�g��ᑱ:J��H�ǉs��q�)�G1��ǎG�S�Z�'��H����#ݑ#��}bxN�|=L��B��kn�'LC�����l���j��%a�Un1X�frkz-.�	g��*��ܵX!�JF�"cmj�J���~='��[<1�Y�Z����Gc���t�z#�n���W�Q:4�'n�D�-�:���bJt��<TU�a�X��W|�?>NvD�r#6�0��0��NJ��b����RKq���WW�6��1cSǏ ����'��R�uFj���i�9���M&x��8Ac���m�_۟��{o�k�F|-=��&w�G�MཱིM�E��^P��t7fPϷ���RN!�.D��C>Y
�d��F~od���5��F K#�V��I�^Q6a<sS1L��ҝ���;����~�"�BOL�Pُ������p9Vj �܆��M�G]_�� t&���� �6gi2:$z�8���xL���3*�qok+�W*﶑�Kw+RNA�R����	��ڬu���X+�*��c���
 W|et��?�r���zSs'�r�F*�hC�u��jYc�Y������Կ� ���/�yRM1D�S e����t"��s��0>�0K�ɳDH��5� ZS*zˤ��.��� mL]ɅvV��Ol�5���Jc�ء2������#quQ�q�Kg�ş���E?CC�:4��"@�R�����7��YC����z����l�D�:�k��#�R�k)"P\���IO��T����n���[��;;�8+Y�1��%Z��TȺ�U����J�&㍫Q�y�2�ι��Y�2s?	CX&����~��y�45����ũ��de�����eZ�'�F\C��(�w1���sH�e�'P�c�C$�Q��]L�ْ���bl;�MeG[�c�؅�ޚ}����LcWW�� �������a�3c$�9�8�n��
6aJb����ԁ�]�B�� z+,�TK^�B�W�nx���6Dy�����v$A�R�0H�+��2��X85'�
H��'L����'w����$ř�*2�Ȅ_/�H2��6x�=��!yB�,.�k:�F�"�����f��X����oP���:�@I�q����%
��������� Q�Y�5� ��~��G�A�˗�r{��C��DS��i��v�'l=+��N�k���[����^F�Vdi��6�<X�Z2F/H�`Z�e�.t������D�G��"���v�dY�<�I��o&b�Ύ,���7u�r���vc�L��r���`��z+��?B}����|#�R��<f��f�a�{߶\6��~C3��]�2�����|�fd�p8��Rf�k���=���$��,���
���*��ZQ?���������	�M+���uZ}���27��f% �Ǭ)of��/��;��4��~n�&a?'�"-�B?01�E�[�;���  `�>�;V
�Uܯt��9d3l�}����.>S�|�%Jwd�{����ŏ��PPG���8��S�Q�6,�3i�VI������jQ����t�^,}!Vj�C����(��	@��@G�9�֙WOb�.(�&�XH�U�4�=�Ri�I7����Rw�xxz�;BW.��/�d�Fn�RJ���D�#GŶ��8i��8����T�1IH{��7���Cp�CH!��^��;�&G���_��[��{��au}3r������TP~�s�r�)���I�W2��%����D�O\>�W��']W��"�0N"6T������v8<j
��:��Q�+�����fd�(bɉ���%IRJ�u&���i��`8�'�9Q�Qo���
�Yh���߷w������+�?�4�P�k8})������ՖNq�e�3���X�?8�?�!�{I�
��rq���|)�VW�����D������m?0��Ś����ϑ�,f\F
�&�n���&�&ޞy���H��uN&���E,6�������g���Yp��C���:�z��&�v�ߗ�c�P�4��O��Ps�����iN	��p�����>�2����K�+�&�#����cРB�-+�4M�q\��SJ�����M��S�X)[�`���~�ڭ!�q.��b�w�\��v� "I+&Gk��a<���mnF/�&��`��Tן�+�����&�M�%��|�S�#�.k��6��b��>-���cgs�P��`��˯t}`�D��>��;��k�q��r�k���Ԉϗ)�d�C!�-Dnr��p�UFNI�Q�r����a����QP�4΀��|U0�F�������W�� y�@�ɸ��`Ӳ�m���z�]�:djr�R0:�?�7���v#1a� TNQ�FCN�� �G0�D$*�2R�7"W��&H�"��	�8C"#ȏ}"��ȴ�lr�$�5>�ҩ�R�퍁�[%�VdvT$�K<�Z�a�'�x,�nWbn���a�go�9��jC��TI���E�K��?2}J ��aO��sҽ�܀,(��667��@2 �!��QNn�]`9V��t��?#G;���{<���������r�)̍���7OE��f��/��h9�G�r�~��Ik���QM��5E%��1SKhq�[\b��f+��T}����^�Y���n��"�o�/��3b��y>�`����`W���p	�\T>eo�Ɏ6vxl
��߂�n4���(�-ެ�-��٥X	j'R�TX����:�zp]\�\נ�{��56#��H�4l���:l�5�����~�i� ��&�=�S{7���~���-LM���z�-n	���Kw��mJ��Z�<���>8&����6�"a������dM�f'O���M���γ��|�t\��P.�����>n���&��������pI�|�Ҭ��a������T�"�����\)�H�|��q36Y�,(��g��9����0Y��7����/�t5��%�d�)���v2�ʬ�\��Iގu��;$�8=S�}�"7�݀�,�U���KP�J��&��L�+�b?r��QX�ln��A+��V>n�^�n�4�O��,��r�q]	]�ƈb�O���hMs�m�~���m����J�OB5%�mU���P� t��'�
Ja�#�9?L7?v'��z�oId5�¸w���V�:�TޕC�g�L��,�����Q�m���ٙ�s����O����ּ�H�0�@t�x�	��@�뚌�eU�Ȑ�P��l��#)���ؖ2��L�/4�؊�n�X������_�G�ħ�%�73��-��𰊞��;�3��rd��$�?3�%�-�O+��I��"�fv��1pN;�UW%�[�A����P⫲�D��Ry��x������T�}{pn��b _}JQ{y	P1Q�j�P~� ��`�������l��[�q����\w9s吷�뱊��P�\9�����&��6�[9�u�f���r媼���M�F�gd��0�i�^�~G=c�x�	0f�b`.%ri��<W��W�}:阪O�C �_V�CO���S����gZ���Z)y�m& 5Di% �]7�u����N�
�0�\�>���D��=(O�H3�
Llx�W����Cݙ+s�OE��f�MFS����I��߽�L�M�20$P�3ٳ�����!#4E�A-�I�m��Q��C�D�m���V�-2����"i�z�_�����GW�>FWUq�
�q�G��JC���oٰJ�HqI��N����	5���	ֽ�"�������ǂ&���j;�- �ro��RmeZ�j��~yk��,KO���&#�š�aY���C;/�u�J��**6��U��ck	�B{���fտC�u�Ůs$8���oc�`��[6�c`�v'MMi�K�k�u�׊�&Q��P�T��|lh��+F+Y`�|�2F���w�+��t
�TA�uf�L~_o&Ͻo��	a�.|���s�>/�⭺vG�B,� ���+�y�8ǜ�G���-�O+zwX8��V�,M�\K�<�u*a~F��&,���1�?�	����y�g�ȶȶd!��I�����Mx.ڊ��fc�Y�{�A��?Q���́�R�Ҵ67�:R���+N�ǉ�U)iQ����A�,�ӃE*"��aCy6�<�%ϳ��������vŧ��<S6��Z�v_c�9���Ť��s���|g{I���
R��*�u�}��� 5��#�h��~f��6�lAP��ن�ё��%�b�#g�G��q#n/�R�h�DwCBy��Ã���Vs=As��#�w����-I"tdځ��xY�����`�Jv�xeDdA��
$��?��:�n�!P�N��ڦC��0��Κ3� ��$+2D�t�.� ��"�c�L*������AC�wkp�A�z0eSlj˧$Mp׺�68ԛ��ӔU�_�;�1c�o���6�"�0f�嬩``�JQ����槪���dΫ���j5zC
Lkc���w,�k�"l��ȖX�/,I-�_� �����-�{�
D��!SK? �c��g��v��#�%S�:-�t�����
ޚ ����"��T�Bگ���F$ �os��IlM��O��8u�������*z�I;�5 ������9��;�תK�Dq�L� ����}_�Y���x���6�, r�Z)�z��<Fu��*�e�o�" ��L�J%n�&x[���oy��;հ�eՖ_`��Ƃ�$}X�88�(e��G�wn��3���j|��L�F	u�/[B���|��ԡH��\I�I��0#ƶ�32��U(|�ɗ���+!%�ߨ�D��8�ND�]Ξ���+�N�no��>섙A�)������j}���y`g�1���
t����O���Fr�gk���b�l�GpvA���+�=J�Y�/�_�'��5¢B_��KҊu0r��}g_C��ל
QZ��"��Ր۞����$���p�9�ںI ��?�B�Dm=��X����"ݚ'�n�����m�P��Dᅲs��4L;��rjD����p�'�޺C��pM���aqk��*,�eEj|���ShAcM0�'���^�<��i���6ǰ�ht��m*�&���bB���C��|��`O۬X���g��)�&/�[ ����v��Y�]y!�O��	RI�� ��V~�G�}n(α]X����0D(Wmj;�=���3%����\�&���Z��eSq���C1F.*��Ev��w����-NkH;�	"�$C��lQP�g&���;Q$��*qŎt��Ƚ�s����\E-{� x�@�s���1�P��n�sTt'�B�����A����%*&P��l���1ڑ][��]~��z�rj*ДM�X��r����j������b_Qb�7�a��,��W���B�S��Y�.;V������i~���2���o�d2�Y���9��[+�B��/�^L-�I2�5����;fd�/����-Έ�_��@c��Ml�>�`�j�~���k�ApG�^�]�R\��P`ǎ[�;����ԝ>�4ơ�ɍu5�Op�qL<� _= �Z��a������D� j���%BQ��Bxz��p�k�;�}i
��� �x���y., �ߠ��>Ď,9�]��1�%���Lno��\踯F�����^���S��#G�8���%�1�>��VD'�N��Yp���cf��'s;j}�r�S��J+Ӥ�&�b�sw	�L�Jh&}�Y��C��A��i�>%k�B�{��y�8m`��)�hf<��k�?aZ�(�Vү{�>71�(�i�c*�����B�L����z�i!=��lE+͞�N�l���iy�	��,p��%������.렊�/���li��5FEkq�߫�1М','�H	!�u��x�|�7
N���P�p�捫c@P�s83�EP_G���M Ό~��E�u�A�g7�g�5D4��Ѿ�
UV�,W� ���^���^U��D5/P�*��0�Iׅj�df��˿�Wo�h���%�L3�
8D�g���W�AfF������o��HgR�v���Sy�h��$�X��h_�w��k7g����X��o���m_�'�/m@;@�����<0�ɛ�abY) �.��D�^�|vIO��ᔖI�P��+��y�@fF�Q��������R ���Z�ãI�X��Ԯ�n���2�zΈ�3�b� ����s�w���&��Y�Y+K�|�_��Q�Ϸj�n/����5�x��TR�dQ��Q�A\�7��XV��B�gn�\͈�	м�XQ�:I���8a��1�NQ_����Xub��M���hqcA�� ml5a��6$�ʩ��<Q��:��;�zy��j�=�U�h������-�Z���Wi�z�v�T7�꣜��[!�җ�侈T�8@05*�����]��W4	O4�ØMM* �QNb�(ժ�M�3M�@@A8M,�h��Fɥz��������v[�ƽ���o�!c~d�I��Cz�h�n7x��J��d�T���#��^a���6�bï��r�T��-�Z���_���Mu������Q@�E�kb�<{��҃h���u����A=���V8#��6EY�v{F�%�8�Zx���㾎�q��d�Q�X#��������>�?��*���ݔx)�l�+�	it�6(�A��	Fo}>��S}��F13�����*��T\�G����A�� �q���4H��k���E3��{!��5��om�>l��%�S9���4��ho�ڼ�k��?�˧�>�*�>+���A�l���93���1�ݨ�q�/[mN�[)�Q����|����	�Br���A�l�O$� s�p�<�~��Q��f�pO���9v�s�NV,
��-���L����0����o�5c��y�k�A;��!׶���m���jð�h����i �����D��C���M����efl���eN�Cn���г�K.%�ʃ����g��6�7|5]��O���t���)��3�?(���H:��ٔ�ڮ��Q�Bti�yǃ�y�`�$(��X�m�?FR�ܠ#b56Q��>&��`�4g%3_�������"�y7���K
%~auG�<��CA��fe�9��*���qc���n|X��-.|�/���g�ܿ0�/QJ$-�U_�D窱b6 �RE�>}FH.�y&<��wxW]��/�{�g�(��;`�EX���igAN�Ѥ�2Ƹ���;�K�魝u)��N�zѱ��|y�O��ެ��M�˻���m�����Tgh^�â����3vו�j��O' �o��#Iy7�,=��G��3�����B�U���<��I���k�;,K�T!|�#�"n���2�T٫�J����%�V7c\>D��셓��tWyV@�4IJ��'԰\�1�x𷥊�ڡ�<�ۓ�Ȱ;9\����[HDi��\��D/fҤtg ����(Ε3/P�3Q�.4q����g���j�X��`�	
���Bk�:�bR�5�X9pB9�gP%�B{`Q������)�)�p�	�tV���x���L��n�c�R8�+�ӓ��_��B(���[���Z�q���F�
d�VA�P���l,����J�>&&B#Q��t����������.�j�*?���(�AH�:z@;1o��ڽ�'ڠ�%��Ԡ�`�O�ى(��g'�5j9�.��G��d7�Q��� ��K�S ��2p�'Z�}��l�ߓܓ�2>�D��\��K ���sH	G��.����5�����`J���y�n?��.B�Q
X�ÏO\�A#P�k�3\!鼺��g�R�E�/�r�A�� 
��nt+ᕆ��e�oy��I�ʽ!{6�?��AC����_:5��U��N���b�A߼KY<�B�l�N-'�8f�	9I�7۬����s9J��p#�%�	߶(���"o��5�W����^������R�s���F�3HS�!N�َ��(�
�K,�ʐ�Tn[���T�t߽�q�����w��~>KC؟YA�ln�<���-�So��w�=�=���������Zsu`�W��Y6�W����:���]OH�ߗp�R>��� Օ8$����Z#Bh+��LLvDBE(�V٪��xV5�"�����4�y����[�1e���҅�2�z�j%�ژn9��Z��3��U�b�����ͅ�/�����Fqd�ȸ}�_�D����c%qE�E�,܏|Sw�г��I�-ջ���T>yW�If�����w�Rc�1�'��;[�{Z*`��Ⱦ�$8f��{������O��]bX��{����>��54ؗ�|�s����E�7����R�A���-�(3�%�Ĭ!|BwZ'��Q<���!�G�/ i���L&߼b��'.(FDͻ_߯��c� ���܅8��7u��z��J��ß�5��o6�)�|�Ǔ�l��R]ٻ2�2=�X6~���X�b�Ik�����u"�c��P*!����R+�y�`&�I�9��e=����aQ�\r�7~�"����s�b(���	}*���H�J��q��i�)W�)�ނ�D�/��9�et�VP��weI�x�)�3Z���^�*���zu�P��x����o\gt���:)5��xi���>�Lk�v���Kux��6]%���/�"�r댴�J ����{7�q�J/̠�tm�����׵�4-YH��R���N�㍭/�����g	OG�)�W�{��	�F�O��ʻf���y���	 ����G����)(�	L�P?���V�.j�4I\9HZ?�-y�5آ��{�q��ԹCyB�;`IT��R����؋�˞��pY��Ӛ[!0X��I߿�������3>v��5oJY�� ���KH�@��\�ɇj4�D�)^g"w92��a\�R��
�qý��|2���bt��Ajwiõ��C��Z
x��ga�������� �k\��ooE��C����BkLl�䁄�d�h0�~f�/�"#�M�˦ڦ�oh~��Fl�+�����۔ܑf�@�����mH�n�~Dۜ�6~�Xb� Ѝ��i}!��Bb��(W��ɐ��hp������#;����5H��.^ԝoO��k�Vb��}��������1N���3w�qM5��?����v�"��I� C�y�������F��:�>�>��-f�Nct��:+"wA��� ;TlYL 1�}l���x��IW���
D��{�"���J�ݖP�iX��Ho\wV�r?�� ���"��?�	���{�� r����D0�&<�R�����YW�s�$����DV��*N����m���q�F��7tT4���k�c��t\��X��B8Ta����[g&/V���OqQXv@W���ޢ׉��c�gs�B�&`����q��d�{��S`ڥX>�%��Y�Q���5Df���m�d��JhP�Ϛ�A�I9.^PM	5��^AC�:Y�gHv7�7;�������T?$�Mf�ܔ����_J�v1��
!��:�A�	�X��F|�p��凙˷��^5��{�<��]��c$����hhgѕB7�ܰBD�e��Hv쑎Ѿ��	,ޥ�O
�B����:����� ��Hn&N6����Oe6�	�y~�+<��L���*	T���J�G�"�X���<0��2Hڻrhӷ�\Q>���xO�j\�^��Hx|V�����֦C.���ޟf~��X���4k���Q�.Bw+�!-��. -64��H 1kѦw�~҃ul�����q��Y4c�zX�8Ꮾ,DBl�M���=rYß���H���(�ue�D�A�C�{Ib���2ҌH��Y��mg�����LRZY
f��-₝��ԟ����RK�K1�m�ӴMξo� ��������vϼD��D�T�=��8�������r̞���0F��zj�Y6.�,�kkx����q�(�	�F��mh�q��WJ�$�ˇ "Ɔj���G�NLeaSl8�^��J#��-%#�`w"7XZ���M�q���
�"=D[f����'���209��Q��8���z�ב���w�%�I
�oZTo=���B���*=#��~
yHt�Te=c�%hW
��%n��G��>̀�w-�g�E4��+nz��U����juP�`�C������%{&$ Z��x��"|��,�1b�oZ4Wk{A�]��Q���ok^o���2�z�B���2�)�ʜ���(�ĢD�7�i��<��z���,����1��VTR���z��Zf~���S������q���A�p5��^�U{˪낒��Ek�]F�D�i�LiN�s��98��	�ڎ�|Q�I���b�fJK�>�^�A���҂��҄��Z�&s,��D�DĴ��|<N� ����W�]���G�h�O��ʥ|�ZH�7��~��+����7��4��/$YU|�*�Q=��)C�������8�݌q;����n�u�8���7���a�\7�`qN�>F���s��<�P&�V�0w��col๖��dW�B��#�����z�la�cd��$x��x�b�e���̔����!�6G�����SmlUX���>Q�*A�s5Mk�,�B�0�t G��S�#}/0S)u` |��$�1GLU�Au�������%�7�7Ni7����Z��q�أ��]#B7�R�٣��a����e,Б4r2A�^R� &G�l�P흿�Ā�5�ض��ʆ�RW�`sA�S��k�k�:�z$�~Xؔ��W�����'sܳ��$%���4P-�\ɈM���Nl���V��V}� ���_���a��LQ,9�|Z��*�u'�Zo:�7r�E
�?5�Xee8��������o�{|���G��Ep�@�5�?�x� D-5d��kE^E���Q��څ �����6��#x���r�+�=|�c#ګh}���*4���+��rK*�lbY��p�ٛM{�!7[;E�Ҷɾ9.(�Zn��.T�����~��E��4f����Q���q*�#�A�̄ܒ-s_�xk�P�;���RKm?�c��a����}�+
�"�+:��l/����~�֖֗ې@ߠ�/�q���N�^\����9W�L�C���C�ћ�EB�ƫ�:�t��X��-H���X��څ�W�^TU�6�X�K�����y6[I���j)Vg�=�藾�����r�	��l����T�n�-D�u��v�d����E~)�l�+[i9-%�7������zqd�����
m�~a���:�SkQ�@W�j��x:Q�@��(3���M5s]�����IU�v>JZI
;W��#�Ȗ~��S��~��?
��w�l�4ǀ�������K�LA��&�M���� �$B���c��Ã��/�9+t��r͵X�J�gK�ْ�]��X����j@șF���l��eb�����K��1�0��9��j��f��RCc��"�a.��b�� �6NZ��U�u4�I����Z �Z߯dZV��\����w`��d�r�@R.�RG.��iS�9L8�2�k2��Q�X`1��w�2ue g6`�eC�T=L!(%}
YQ;��O�m_ף��O{�)�.��/�hfE&ĕۦg�l\<�XgN��$��,m�e�J�<�d�a7|R�A������OD��`w8m�h�'qU݈�A2Cq�U����Ŝ�Û�����r�Ɯ�:�����\�ӞA>ߠK�l�qw)��UY��h�����/cZ?Zٝ�����Y�^�4�\��b�;zJ
�A�%����s9ܗ�SX4w0��h���86�m_�����b^�%�q�8�W��-�U���`v���oK�f����lV��ær���:dK8�"	�?�a�����2��srD]>���n�-}4�p����o��W�3�T�"�pŖ�d'�)K�e�g����F����d{
�Qd��̉ߏ���
�/� ʡ/��1�Q��%4jL�� �d�:��J7`��Ռ.�������XQ$7����nhG�c��_5��=��,��]GPь-󹃳 +�ͬ���D0DϦ�}��8�]	�_D��Il�ˑ1����{ݺ��Ĩ�~�{���[�@����a*	�H�6�ȼ*�����8~���m�5��G��6��,��P=�1��s�1����M-}�i*渖LZ����F���񣆄�.U1IG�,�AP^x���/~�f�������E�l�\u����BҨ~��s`��]�0yM d9��<�<?�i����`�W�_��F���7��I�j�_�VY��,�J;W}xc!OHԎ�x4���k�40roPŬ�W=�C�,�ę�t���}��ƹ��{o��H>�0�Rwԗ���}MBW���-��M���lM�`!V�&b��������4�(a�9l �Nt[D��A��J:�Sd��`�󩕡�L��Y�%)[5�ǖ�PL�����SӘu��)P}�Qۆ+U���G���e�\j/@~ˠB��_d?�@x$�1��S7�#7nV-K���G�Ǥ1IТp���i�/�9y�y��ě<Z�M�N�qZ�L��d�9daj�/Bp�[5g7\�F�"�P0Hq4���(J��㛠�Á���i�w��/���~Qk_7&|+%���i�	,�T��� ���~0%��۞����J4�bK@n�]��ٙ��_6�kE�:���s���s\�2P���K%�V'�~����n>��)'q�6�`B�+P�(9�P!��'�C=�?ݩi�+�dWL�LUkJNR7�Y�Y�T>������I%�����a��.���)�02��#�S{�̃Oh&Aiv`��?����Z�,�Pw���M���A��̯A�n��4$�jI��΃��it3Z��^�c��|�t��(T}2|S�2H�ۧ|�����9K,]4����@,.Z��c�u���&���e�����C��_/�%�}�$�̓�6N�Q��b�]j3p���8�#�U�Q���V���G8s�����/�� y鐂ݚ-����-D5x#ܤ|,Y�Z
�!g` �����}��Z�:3�n�s^T��Kֽ_�y�M�XR�v���P�qB�G7�c�%�>�!���Ɔj�`5+�bx��%���[q��$ŗ^&aa�`�r�����+'ߪ�;/�K
���z �K%7TK~��}"�ɤ1kY�㵋t�#K|���4�;��ʐ֘�0q�'+\��[G"+CX��փ�7�"k�c�"6��L>��B�saB��;��2w>������W��ܓ��v����/�`��U���&��e��ǅ�G�{��	E��<�0ܜ��s�lK�v�+D	.�����O<���R���C�+ޗ����j2�i��l�ŉ�	aּ�9"n^��\��s�c�˹T��#��0(�h�.o��'}q���y��^W�f�d�x�'�uMݕ����ͣ[=R��	���OE�9��~���t(t_.��F����|zp��T�In&8,"ـ��Zg�n��ē$P����E��j�Dg�ӡ�����<�@b��g�K���{�ǺjH�������g��N�^Pl�8��i�0�"_��D��7�s�(hԼ>㔭����G�Ȉl���7�ŝ���h��l��(.B���]Ǣl2�1�O�3�N��z+����U�=�dQ e��p]+��cH�?�T�'.�U�B{�״34:,��vѶ6�.�é�ͽ�SdT&�Hxܲ��:c� "�
�=TB�����W%�(�k��Y' Z�w|Ƽ�E(��g��ӛ�S8�.�p��#̠JJ�*t u��3�~���	>&�L\�#F��a?J\Y��sK����PG�	������w�b�:�l��[ZҮ�@��yYqf�,mD:��!�������:�))��!Z>k&c.�:F#���16P8�=Ne�����Ȓ����Z_�3�%�\ܑnE�<�}����ɺ���{��-���5�ѐ$��<
\j>�c������z?E���e���H��I�X��K+��C1s�u�l�9�Tp�}�k�Y���c�Ѵ�Լ0�[�9n>�	C�]�W�"��8}���Q��F1�_�O��B��vy�(��h�	���gȵ,^��$R5C>�;��F��DJa��Q?;P���I,��6��b��Q{y�v@u��A��6��]8�!��w��򰋪H���c��	�'2`�W���Y��}�Yv�P�!����{Ca:.�§�^��Q
bIf��G�<�qO��:&�53�_%3��[�%���Gyڮ�I��M��ɫE/h�b�1@��;7����.r���0u�0AV��'P�|yf-ڬ�*~��a���)Ϗ�uSx�%�'���Z2�Q��~kX(�X�M��\�m�P��z�����{��ղ����{��>�Ш��mS�P�BmFaT��<���0'���[4��%>"��g�1y|n� ��6Ʈ��o��q�zѓF� ���7Jt���^ɀ�Љ���4�$���oul@E兜�_4�w�.�	�X����[��#��Ԇ�\E��Bkxv��e2}"��g}V�\�C||:^�]��=�{$�O/�ֵ^)���8K�"Ūq>.��h�@mt�-�[�j���J$�����Y
���s����293y��+���p98h��$�УQ{����{>M��H]0��qB�=i����V�`S�K���^;!X.�]�H/�tN3�Q��������{c�Ի|;/l&s�a/%m��7y��3_��ت6��m���њR5���Au�d���X��2q��ܱ�\7P���y�i�.W�{�ja�]:�b�304�mV�&�F���ȏ)/�횠�۽ǁ�9�l%�ZM�r{����K<w3���Gz��hc�]3�N@���e�Qw��Þ"F���R`ᇘ � ����s�����͈e�@Im�`���l?�iH�x�C��#1��w�A��	�.�0j˸��Ȭ�`���&�3B�"�1��i�F|��e�8�K6����w�5*^"��ӿt�3�d)`� )݅�i~��hCg�۵����X����Z��q�$^�Dյ�G�����z~�T��Jl�ѱ�w�~#��O��t�&}�V��;�},�����b��:ӭNp`����(�`g���
,'�8]�`�qn]�b{
��&4�Q�4�5�:��A�s���+���F�jC����	�ԚH�F62v�֓ژ/p���'�*z��,1�UC�U�����,�4͌���B�m�Ef��"�,��Q�'
�[a����`e�E ����~��I�_��& ��B��wЦ&�=I�x�,G�Uo���ua��Q7�a���+̠"���A߈����	Nq�X��h�w����!4k��|-�}�/��ax6�r�[Sו�8�9�e�-Օ�	8>=N �U��E?w�w\<�t�f���a�S$+�V^��Š\[���	�˃�Ki�t�\�ݾ��+K}�dV�a�#��cT�ܝ���o�	��I�-�I?������3AE��A�O������	�к�Z��6��RxNdV%|r�|�1P7����yB�0L�/� kCQ�����V+�y�i�P�f�E?�EFǵ���ū�X��*��i��h�ċS��e�=���+����)���hژ���Ƶy�1(Q�����\�꼑�8�^1�ʓb�u���w����G�q1�:�Qj R_�[DM��r��T锷��>61��k���w�7~`�+�a-���M���?�T]�6�wkt�>�PR����ɴ��z��x�l�W�0�bJ�kO �[+�N�llZ5���3~��!G%ʧ��w��&�L�,7m�'��'����4�Z�v��I��G��_�5�~ujk����很�ѱ+�1��D�<�wQ�!f.�4���H3(v�a��-o96�Gx'��+k�?_��5������'H���L�b�>�Cv�#sO��g����A�]��2�~O6�[w�{�G��*r�_U�Q�iXZ����eR&L®8(���u^�����ԇƝ��F��|���z(Ky����Z�e��i��{��vZ��&��lX?�i�#:����������bA��0W����n&���Ω���;b'�nT���k�:�o�ME�� � s&�q�S ��bZ[�t�M^x�9�;��pM������s$}��:g��a&1N�1(�[�C"����_�BS���}��N�A�f�_R�~�Ŀ�Z@<Wj���e)�:7{�*H�Z1��6J�Zϐ�;G-|�0��Q��@H��Gpp�rp��"$h��.��g��6?r�U��dܼ^f��'�@̕���B��g}!���|jN��e��L���poC�����7�� � ���H��,��Ã�(������i�Z���Rs�?���Hq^�(ք�.�M�ͯʝܮ�+���gq����5���>��R�5��U�VE����H����V�f9Xr�^{׃n=?����A8B�V��j,�@3f� ���t�8�VpVT���W�2����z����̓�״��On�[�V�-h�[y8����Y��2�گ�L{>��Ay��(Y�(d�^�
Q�_Q�v�r� �E��N�l��js�Kx'}�Zr[������[���&K�Щ��a�{��a�H��[A�\�&l���ʁ�춰X�е�.Z1���'�!
5�&���Ò�B�qu$�z�A%��檉Ha+A^�ө�s��D��n ���N-d`�'�� XUPo>]��߂��	!�1�r��B�$�@���9?U��G���:�
���uQ����&��K�C׎>���!1��&��q<px�����`N�F� �������Xi^<���q�Ra����ؒ��m�:y&��u*�p#��L���sy]�}d�?�p�Z��a�.#�Y��Fri��ߵ�W>�pP��S�G�;k(�`��_
/H4���/� �G�]�3��A��i����D��ػ�y���r��rv�̴U*3y�qt$��x��SE�� 4� �V�чHx��$`�����%UA-^{��c�_R�����Nhe�_�ã!���Z����/��k�ԷD�[��d���ԅ�l���qAh��/H�������s�ɛ�#vk�κ�O���8��������SFp��3���C��e�\�)�E�7��l%R夊���y��s� �m*��x}#�[���~o1�{x-βj3K�J��������h��ꁖ҇����Io�b��í�ȶѡ�&�����E�]�9_��1����v4�)�`53�Le�"@�0��)��'^$ii�� -y���JA�#̿N�u�L�T�IO����������Vb����-n4a�'��!ʯ�PoRƋ<�3�p�uw,0��v��2����y�:��Z��_��/��\�ƠFq�_�n���FU�H��@vҙ2�]��0+�[Q��0�"��
�/�7�$X>�f�v+ww��ϕ۶�����˙F0�O�=)���h�#ʭr�9Dƒ+�_R��Wy<�!�m<ع�g��:4��â�=�nt����÷��r�֭,�6BR]�	�����5�eM����"�u~&;llil���Vi4��e��z�1�7���R�D���N&�ȇ3Z窛�ܒ���o�A�i�^#��D����K�.8�){&k	B;h�0�]-�@f��"�|E��Im±��9��1��E{���R�a#�����M��N�ۢ%��'�a��ӱ�!��h#��ua�eT�.�r�L����y���C����9���B������
2ִ�J��Js�D8�6XMȞ���՗ҞpfC���Ǉ��F#jś>�bԿ��/���^ߧ�q�3�k�x����ϕ<7־ĳ�"VF�Y-q��B�)�s�f��~�+Z���I]O ���6\���3y�P���s�w=�ԍA� ;�0c��K�M#�"���bNF�KQ�z���r|��壖
��yK�֥z	v0�]�����r"�}��K�(T_���9$e[.}I%ԛu7�����둄t�!�D	.�5��a�����]k$rt�j�iտ��1�rN8���W�xI��S���I%״"������Q��s��%��r��3��竘����bUSN:��e ������z�h�#�J:�H,7�E�h��,�;��~���^s��A*�[I;'���z��1#i�sX�x?��ՏȄE�/������!j�ұoа]`�vx0q�e�)����PeO�=�A�dGo��e.�i} �}34�����d@����@cު�'U.z s��\ub�r��)�E���7K:7���V*ĈV�4C���FI���$��BgO�LN��|�U"�������y"'�|ذ�<}�8�:/��G�(��̬�[�$@��&��3�3�~�5�!��c*!}{�a2��2{���g_����W,�y<�"�W�m���=,�;,f0'�����(�ꢼW�����O� �:�3T��<����&%_�
Dl�T�$rG����\�h!	Z2?,Ee�Ez�&0�>Lc�]i:c?�G�_;�l��ul�ʺ1����J����I��P�uOX���z�c�.�WvDq����d���Q���S� ��@�M����M����C���ݢ�x�/�@F��_�Γ�����+�*_/�@;�@-����G-����%��vI�����d�_9�]��`����s�ʤ��$׍*����ZѬ�73����tKz[18�����Xʲ-�qa��Z'L�g��i�/�S��/廗��5QA� ȘD������T�ex�m�	���J�=�ls_!@��fE���
'���MDL�|�����Py˄���Uw��&��l�_�G���5�;[���2yB�A�i�*=�e�� ��
�Z=X*<�?K#��� ��nll˩��W�T�k�'�WY~�l1�t�|ʀ��4��r�����=W��&�����Rd����c$[�s�y��;���5Y�U�yB���s�h9��B��3[w� �3U�9l7Z��H�}��� f����x��XJ��^��+k)����NLۛ�<���4G�<x��c`c�X�Y`�/��o�V�R\�]&����
��'�/�"�9�t:,�
�6w�Fi�����Y�܁�\~/v��t���:�C)wUcƳ�1�"�v��"�6��=EX1�V��^n���~��nvP��d����W�7�o��,LԳ��F���ٳF�o�Rw�;\u(��.e��6��+؎��P�y���@���z�D�Ox�i�̰������lp�W�i˷iʀ��;��*8���Xr{�=P])u�_W��|��x��M>�>�+�͵�f�ag>�s�E���B��*{�KSlT��w��^�4f�l�*�c������il�F,�SaVH�����������O���F���������`2�Cu���b�de����8an����\�$bb�{׉7ч#�{���+�,p�m����Xd�Z��VVB����N�j�C�`�2���_�e�LZ����9cL&���1Q���,��/ŵ\À�Tя/J���/�1#z�4v�K:��~���8p��x7�Ka�6�=g�7��k8o
�^;LntF�i�DD�Nb�SB(�F��h:,�*`���ƭ�.��e�N܋�E��
��
�%l�ZZ�=��.��ܚ5�t˅��"�q��7z�Xʗ:����3����:����'�<�\���M��hƮ������p(��z]z��
�ש���K�ɖk�1�\���!�ץ��̫��y8��`tbN��l�7����c�o�U�[s�[2��0(alL ��@66&��R	Q:��@�����\#y	�뛿�&�[}���)
��?��;4�IHN�X���w�4��]���N��D-��8�Б�_��4�,%�g>��r	S�1a�����ߖ0ə�W� �q�"7RI	��G�{ݝAj!O�L�9�9��e��t���s�c'ۡ���lƞ��P����*T��+�8E`"��cX���8�'�[UN�3oS�M]X5J`��!�q~�Y�S֬��Wf�s���Y��$��_xIY�pY�+�u��|��Ѫ�D`�y�m�<�Y�5Q�7�M��� =��^�=�-eS��K�dȀ�n���8�V�Lb�y�ۑ3�2iZ��j1�Cx������'h�>	�����L�yGs���?зq]ȳ6+r���E�ۮNLR;/����2Jd�4Iv\'���H?9���<�b�4kqml�1��gb�{�����.�t��T���tW۰�)�y����r�.���B�ź��@���.������ڨ�T2 ��'�N��jF�n�����X��J8ŗ	��gE`!�&2�+]���p��}m&�I�mM=m�J+��� {s�:�[8Z?T�k�ᖚVf��k��)�[SM4nN{t�猍�v{*g*Y��Wuɨ���m�3���Ʃ*��!��RjR�����g�L�������SБ���޾-�%@�Wp�=��]v�ȑ~�0���A�A6t5��+�lLG��x��E����[S0���[:��Ն9>ɱ5tP���|r�L���5��4<��\)��#���r͜��>&M�5FYaJ]��M�u�߲L*#���W��i�2���|lW��Bh!*�'���� N��1X�-��0�+B���/��Q�[�����-K�[\��t��}��^x�ؑ�t'�X�-�J?˥�!����\���Ki=����G���̐��\����>N�����Lz�ݳ!2�����R����Gt#�^� ��4����8~�Žb�c��&���k��B�P�[�H�k3��^�����v��vd�X��iҕ(q'�V��H��	b���ޒ�+�\�8�%{�a��*�-���w�1)Hp~O��Wm'"=�:���Y�J�pi���эܓ�¹��|[���,��wKEWݦ�����>�	�","�U^�&���ٴ_���k���d�P� T���/��q#�,��,����Ў��{4:���>�����ޚ�Pe�g�G�m�i�CjɈɋ�۟��qA�IY�,"��H�<I��Lۚ5�-毢F��"n'(cބ�� �W��u��_W��|�E�h���P�'^Aq3��A��r9�P\ڞm�vڦ9#�0���0�|��}�3EY�:L���E?Ж!,��B+��Ks��rfD^�������ه���دs��Z|��2�����,0n�L9;Y�̕��kp�<k��.����M����ʻ�+�E�
���zuj1q!��N:�?�"U� 6�CմVEt�9�Wh.�q+)}?Up�xQ��6���)شp?�?K���9@���¦��A�����g�T�ˇE��G��}r��ԝ�kg��%���Ȅ����8ù`�9���<JV��m >�T�)�n���k��%J �A���H@��S��w�2�D}a�>���[h"���0�9��b���V�4{�pM�k�_\�K�����ߗ�s���^L]��nď�W��Eu����y�A&M���+����D]M��9
�������_e�/�&`��0bG��y����o��=��Jj�q�������u( $~�S�K�d ٫m�]�G�Q"�������Vak W,~�!@�=Гhg�o!H���xQK��F���G�N
����־��ޒ:а9���Qk�5�6D���¼a�8,��c���c��	�7B�^씛�VZ^ylW������4�X�۬t���yu8�&XD*����:2W�Ҕ�Ϟ�7U��[�U�Ɣ^����M��r^�u�i	*�Xr��<�K-ԫ�Խh��~�t���he+�`���Z��P-�S�cP�f����#oĸ�hnr��["�� /�֮zb[��K�%,����cG<����eժ��������S���MG���Fn�e��/��Y��.��n�1��!K��G�	��[�9�&⽴�B6�4����$��6�t5HV�,_�.�����~Y-���ĵ��Z����(��I<;����������$a��Ε���-��Uկn��,��g")xA�B]�<���R�43Rmx�&8U�� ��U+�c�־,���%+��>�Q�t�ý�4i��pY4�ܶ��x�$X�r��ᒎ�[��ꯐ�|d��OJBV���n�:�6�������|[T�?y�Q/�g�)�@�fj���}Ρق�3�|&.����,�/��+x,�)�e��m�n&]�N��Y�~�<ae��ofVq�$�[W�鯻�VjG��^!V��>�!�ޡ�}�d���g7�B���%-�qje:(a������~ϋy��4ϩ��֯ƓKa2��*��|���XCx��4�v%؆�:brޘ��1g��h%��}�m�0�ff���oY_"wG�/���䒆W�c	r�R�8�b�aG�<c)��N�n��g�5��ÿ1�dC�+ڵZ�xN��0`��[G�;7�x�&��1����}`-�Y0�>��%���l�.� ���3.��٦ƥ�$=Y>�vP=� ���&����>�,�r�ֶN��n�?^������3'�����+�uc5�<��� �I)�L3�8w��jC�!3qsC� �
w��M	��b�.<��g�dY�f��~�_r�5�*�U�0��T/��	K�e���)���5� 8܇F��o놕T�P��r ��/p�v~ox���kPmB��l�{�3<i���B����OQp�~�"��Hx��S�G!]'��U��}7�!@c�~���P�Re��J&������r�w��޵(܈�R��w���T�%�?~����5�	�N����ʀ8j^ُ�8�Zq`���f\z��� ߴ��T��Ɲ� `u@>5��m���\ei"�_�.]�BX$Z�H�R;�P�����G�&�?��V��P>`Ƹ��a6�
q`�������/q�c�g���
�v�4���Zw�s�I��XM����w�Oq9����XT�6��|��L�={�/r4��6K��p����S	��*&Wg�2�N�@a� h2�٣P���`U�e��8�)a���+���=V�u���H��x_��ڞ������_D�4C4N{��^�"���C��6Cw$y5ami�_�� P��J�u0C��5!x�l{BD;�i�Ȥ!h I ���c��Nb#Ζ1�/���":�L��O�^3^�uK�u���}����*X��F�rt��1K����z���(���3)��X���_w����Ġ�дK�]e��}�uҤų��n��]*M��=8�zoN�I�n�+�:��E�eN�l����3 łuK{B��ᒋr�IYj6���-*���c}!w��Q���_J�'P���ӥ�_��r���z
�X&�7����D+�J���o��/~���V�iI8���v��sf�8�K&��Z墸�,�,6c�Dv����(W�/��6Px�;�yO.�@�Ҹ�	6)5_k��T�@��O�]�F1�B�5��F3/8��/� G|?[��D\s�r:��Z��
�B��]X��х��w�X�Y�U�F �Vl��T���n�Rl�VE�.�j7��bU�{V{u�(�q-�a�N+
HW�\�6״x�����?�Џ�]����b`:)��Qi˴� Mr|��+�m`�m�$�TC����/WՕ���\-�&D�?>�+"�?*m�ޱ��0��>�����DS1�Fmd��S������r����A���@�<��	��,No���أ�+�nz��!�jg��s`�ti*Vb=t�KV}RW=D"k�@w-��0+旻@��7�@�[IU�9H6M�-B�V�"��=���
t�4�#i��t���Q��]���A5Q�����x2/�Պ"7�\�/5q�Kՠ�B.�_9k L�S@9̖ȇ���敱Kv�f1����f���v��*��b�����k߀9�����\4@'��d�Iv�o�-�'M�+�0`��r�����u;ju��7�}�÷MMS\�|v�W
�
�f�� ��8Kع[�z�s*��N�B$�� ���b��Qk<M!�j�j��HL����F'~}�G��|%���z1�Ì�u/F����v�U_�{�JE#!$.�)��+ơ(Gk?� �[�q�=I�Nn� W��]��HQ��%~c�1�M%��)P��:w .�8�\k�IN��kJ�8��x�!O��N$��C��!V�8?ύ\P�N䟫���p���{��Dq1�c��?.�G�.`��,M�gW��w��䞄f@���፠{�P�=Hl�dD(�# ������#���Y�2��n��$�N!>rD9o���Ţ��2,[_�Z�x*Ɏ�Ӌ_������Җ�:,̤��:0Ӛ�2�t�٨���i��Ib,��C��s���s�9����=��R+44=:]/���T�$ ��py"���|���<ݲ�z��c4�T(��[o3G�,w���58!�m���Pb7%���������b����-1H<�!e��V(QNqd`�C��5"���l�~D}��r6|�Y�k*RЪ���I7c��kb;8 �����Hz���ӟ��<���(cA�aP�TD*�΂6Jw�Y���ɞ�@�)�3[���+�W}:��n��a���z!iV��kXn���D����~1��d�����_x�}q�JZ�.�K�`�Ǿ�\���j)�!u��'*鎡�����ͽ����ڲ�dN%wrV�wU�)&:�z^U,��z�M�b��W�ޒ4�d���J���@�$�$i���b�.��G��0_���o���"����j b���1�K�=(i�x�q���DFz���Ѻ�<`�Y�펷����N���i�m��f��L��Sʙ����n��6iK�{s�%.lu�S	A_�W����9S���^ �O3�>���ռ}u0e7c����Ґ����ʰB��>h����q<��{��b&D�)�1sx�hh�@�}��ۂC���t�x�D�&b��+�(^��?:��{����h9k�������o���4���o��Ҙ��|
{t�� ��`v�_v��?^Y���rL�7����v�A�^em� J}�"H���Q1b�ǍE���wM.9@�s�9�����-Ď)L�}��1Șa����x��"L<�����ṍ��v?u�_�aj�Y�E��S��L�#r|:7<x[߄y��];m
j�	�"ֲD�PG?��a>�N;��f�s�̐dOh���?�4�!N��'U��u\�;���?�I�#�͵gP�Ttk(�Z׶�D9t�ԙ6�@FI7e:֏�G˹w�hۘ �
?B5��W�U�p��� ��3�?#hV)\�]�Y�$l��Iʽ}m%�����
#ǫ��*k���J+��vT�h�p�j���/4�AX����Ǟ��j���gH���&��ᓓ*������U!N^����:0�LA���T��P ~��C먮�M	M�� G�L��{1���w���w�+k�2к	/_YutZ����.4��$9ph�K�J(���2YQ����B�p%�nP���l�d���ZFY#,ܓ�&¤�����I��9Wͥ�0�=yKT��hD@�o�� �`G�w|DJ۽�ˇ,%��?�G�i�U����U�w4[�+���^��
Lժ� �N��2�(�HmMUԓpu2�M���N��9����LL�߶��V�Ao͑��ҭ�C���}j�t,���7�ٙ��p%D5� �/��`�3�q�ő���Ri��0 ��"N[��h�I�@9��XAz0>�Th��R�M�%u�����#X��� �:��
a\��!\��gm5�2Z��<+g^�=V��s�(i2��"u�Α���<{����?�7���령hR@��j�uwG�.�ߔ�#ē�۰;fW!����-j@p�-�)��7*��[�JA]��D��v�V5f2�|ֿ#�%��@�2񮠮K�%oC>��2�Y7d*hcߜ���'X��
���G�;���V��8@�������]����O뭖=\}F�4�//~]��i��Oh�MvM���h�">�+�a}�<�v����XN `����.s��������>�үg�;� ]��8��K9�#C�]%v�߄,o�{zZ��)����O����,�D�쵫V�d!/EV�F���O��o)��(\4[�{0�J� ��C)�����[+���U�D@��YqY~�νv��i��b�P��T��9g HJ�1ņ*�8����i��Щ�	 �y�,�Q̣�E{�]���0�t�MQ�ҘDvEZ��n5���K��zԶ�=�Dq�\�n�C�clW���}UՑ���a\n���g ����]�X+�`
��US�?,\w�컬jB�ܰK��a��R�
[7`F����Q$W��}���je�����@� �Ckp*����,T��q:"l�P`�ē�ϒ�bS���rJ�)/�r�#)F��Ԍ����M�l+���и��!T�xfV.��$��MR_��J!��W!����-�E�mr���黒����E^�J�us�M*���P���{F�������<��m4׶�5�Ui=��7 ���xqy�L�\�l�MXϔm�
�h�Z������y��S�!|�O��)�4�V�B�1������߳h��o�d��d�b��Q�wE�[�2��d��ظ��&�.s3��HX!�6\Cp~XU9����\��r�t�_}��ZK1z�d����'��~x��h����	�{M_�7���h`zsj�a�$�N>D!<���h����ħ��F���
�1?)ӡ+F"�,�O�:6CuPE5۔{X
����
$5E�+ד]�w��J���q4	�EI0�����mvX�6E���'��+�!��;�fU�꧱ݰ�8Ѕ�DrF~��4�v�<�Bf��-�����W������?}Z�8�b��U�6[cQ^�
f�VEI�6�p����7v���XJ0�Y�?aW9o�C[�{�>�/;i�کa��S����iuD>$̱[1i@�G%Ý��]o~O�xO;�i�P��y�������U��gש$�+Rg� {�
G�ּ��	U_0���z%���9��y�ʵ�%��?�l�τሁoʿ�g�����)v��g�d�uvtl,�ƶf�,�)q�:�������㘃��N��q��� Y<��T?1g=0P��v��Ω]A��s&W��e�+C��)�Ѝ'X�����a�8�1��I'j��C��I�G�!j �&��Еu���&����lU�$�}�&{e18+~�|(���>�,�B����3�c�W�t��H[I�h?	9Mx'�6���ؾU���G��F�{RUIȠ�{_vr@�Zo�,�V�r�'������y��eSԑʻ.�WՌ� �����,�@�.��ß�"5]���Dr(�$Wk������aLT�l&�;�*=��_S�Q1 �G>��P���M�Wg�N$��u`wr���\�_�<D���2Y/�YD��b�ߣt���ʇ%�c��Gl��Su�6�#c�q@��.\�|���u�&�H�.m_���Q�0!A�͋�kV��'��'f�[冄���2��	�$���f��m4�5�G60��
�hu�M�;~W�6H�I�vT�>��)j�E�J\��o�3�,�5�
���B_��⢝���;K%A�%^=0�H͛�D��W|g�Uۆ����t^�H<흚)��Z�l���������~��l�s�M���n��E6K4��/#�O����6:�p��Q�����S��V\���عm����;�b�,FOqo���C	˰��:j��@�����&�7�)0^�q���������0Hk�J���G��:����j��x���
��HAcz�]��){��i #����(��!{�kl��ڈ�w��>_���#D����˸�N������0�ҕ�YUh��E�T��׏�M}�>I�1vGԾ���Rձ9����]�z�c���[���'_�?n����M�@���Z�4����B�ב���Z���ҽ�Hc����|�XA�&�y]��X���}�jY�
�?�����16/c��e8��"j*z�ز�����2����Rv�볊qL/��|k�+n"��}���/T
v��T�QQ��1 �}\#UF}��U��$��A�M�p;��d�~����YZſm�(L�M��QhV@�~^����n��:{�S����(��>~`&u� �*x�����>�Ȉ� 5Fô�KGĕA솣١�H'�R�pT͉��Gg����c�o���/|�V�P�3��X�ͯ��"��D��NM�~8v���`��2�oy�ٱ���B%�2cҘ��0�_������/?�X���T�M��zpǿ�H�8����6��o׋�ó����X�w��J���E��2�QB���\+ȫ,!�P&js�_y�ͬu��Q�K�7���qcgӧ�ִ(�;�}ܑ�[���J�� F�J�6���+�_�*!'%���	�
H�}�c5�r�AR^{�;b�����HH�NWAD Hʢ�$L[���L��Fr@_+u�ǯ���c*drx�;���!�Ld�"��Ë��1$U������ϊ#���s<�O���e�hdo��
�8@�c8̄�L��h�uz�T��Ҕ�!��ԩ-�4p=��/!'����_�龽�'�����_-�&u� b+��/�M�b��e�� �ɼj�a�{���6][������agc��=�j�����Z�)�/J�F���Z<|r������Ꞗ�3>���ka��I����_�R�����KgC@�b�R�(�M߳7��C���r�(�TX��039���IT�pF�f�o��+!Q��I�֘ȹ:����8y��n���G�^�[��M1�'m0�,-v�U_.�5<_��bK+ �E���=%0s=���3��^$�*u!�Eې�&���G\bMB��۞�Z�{�;1�#m���Ζa��AV*S�������|ߢ����X����A�V�S))�GA���|��ih���ӎ�Q	���r��w�!iW�I���g��|�S�H!�+zM�8�l�a��-Z��s]�ͦ��7O�Ti;���-]]?
�	� ���!_�9
�v��(��O Kq�|��}�4|���a��l�[<�wC�]`�A���UzT@;�Oڬ�P�9
��n�aGA��A-~ �{T~N!��gF�Ci�x��T�H�`Tr�㶧��bF���a��o �d�w(����}����t���ze^l3�!PLå�D�ُ�ٛ�]�%���u���l 3x�����,�>�O�Hp3?��P�ᜱ�!�Qq+u�ۡ����(T�h���K�|�
`9��1��^�X�ׯ�R��g翡�o����CH�}D��)�S�@���Izm/�C�ќ*#޿lD<V���y11Af|F��5�����y}�kϳS��lD!���s�ĭ�2�S5zO����4����q��� ���N��2?��7r���hm�ͅ��;�q�Obg���O���	/��g�6|�?9�]�;��aL�W��|�Յ
gK��rstK{�iT�X-��p�7�í�B1�'/�+����@KFZ�XR�oG��i$�M��VT��LV�C�u��}��x�	�:����`�9@�n9��%��eqkӁ[*)���;��yi"��?s��2�w��5��ՙ�<ɻ��(ө�;V�N}"Q���m�����c� j���j�����+������!6��)��QC��*��j�QO�65��An;OӐ�#����f�%؃Ix�_Apt����vB��U�$�I/>�ZQ��uV��=��D�}B��_!���T�%�*[EV\�m������ݮ^�u��1��7Ж2��-C��֭�"�0��v�u	�֕y)�֠Cw����R���T>����Rr?�%F��X��g�
F�e>����!�ݠ��s�~.i��ʣ��!.l�/C��1����� "┺ x�@���N&j�1�O,�!�b��/��l�C�v�K��(�i
\zF�om�9?-���փOC~��tt��sQ�	�� �/U]�ݒ&���]*�H� ^��n�'����5�o�����}[&�c�Z,^|6�5�2s��jf��&;?��!W�
�_7C��M�ҋ�!�8���pL���[��vp��#5���;=��u"�IL�<J�UD:Z7��q����D�p���b�D������HU~��}X�l�=���#��Ph���qe���'��V$�������"��H}*o�a|U0���B�,.�܋�Iw�3��m�_4@�KRS)Y+�O?��!�2Te{7t��<��p+j����#��鶬p����n|�mW�מ��05�]�F���5o`��K9���Q˵�&9�OF�5ld9޸1s9��qԅ�HTk�^!�Tajï��)-�qm���^�Yg�4 |��ş[��~`��ی�@�N|��qe� r��7` � ψ���n�b�k�E:�V@=�Z)zA������+���Zp�!?"K�&������=���JY���w U���� 8�}��U���>��4b��K�7�`�`��Z�M\��텲�͐�xW�w+�R��!����T꿡7f?}`T�L�z ���C˰��I��1~�xr�ȴ���DL��l�R(;�K�*��;�B��_�I_���$��ă-�ߛE�g=����|�c�E�>#� �ӒXZ�؜�Eܔ	p�Q���MT�V�&o4��&AH�^}*���:N�
�� X��3��@�i!XT6#*�,D�T�Kbe,T.�`���)�k���"�����"
�m�����Q��l�@���P5�"$��Q�v���y��I�.I}�Q]ġ�\r�6�Q���X9�{+6��Nc 9��p[�u���U��,�F8<�L.e����jd�a)�>!��ڦ����/���,.�Г0F&j\2��O�����rQ�J���4��<�021���>��3����P�t ��i�J i��%C��s���� G��>�<Mz0Oɿ�i�j�kh\k�����9i��O��;0�Ü��Kk$e6�t��7D�5����8J��)����x���M�i�"/I�!sc1n��2��<���N�/��'S�"_ϗμw81�IͣP�_m�D���CL���c�~㟱V�ņ7��҄���κ�K�����T'd  3l��J����E�3��P�h#�V����0p�ǤG�/�_^͵��>���S��G��,r]��ga����j*V|%�!#G�:ڪ��O`2��h�T�7��D�#��X󠘅�)9�Țk��a���B�Nr�1B�KL�0C)U?����F[���=!A�c\@i�6����IW��}�j�J�З8ZYTW�	Y��?a�.[�&W��W@�K4�k�5ٿ��Q5����I\����.QW*nG�!U�)ns3��?;Z��2&���	_;~#jh����}�1L����D;��)��f6\pE�^oNC�V������;��j����(����Xh���a�1�	�{�ʙ��P�3�L���<�5MT���mI��<x�R=0�ڕ�!>��  � ɮ�d�1���*� \��U������-�]{�p�3`)��W]h��x�Q�<#�C�D����-V7���ELT���Z%N�?�vҌ�b7�r\�K�}�A081IM������r�uV �[$��I�'�mf�u	�7łcBC�:�u�_�O?�)F�"�W�cb��0�$� =�ąT�˳����'%���M>>β�@�������Gy�E��9P���:2�g4]������,x��LK֨w2ˤH���"��ej���.�]��(�S5��}l�U���/�|@�y �`� a8���^�;F� �rϿIQ���d�	�����1�qk�"6����H��� ǲ�V�8.lxۗ��]:z�H7y�Y��I��u�H�u$�D����W�_sΑ�-�����,�7 ��Ԑ�n��ж{�6_Z�`i�5F��F:����ga.3��6!�rny�@�=,,~�?�6>e,��2��v�?8LYA�����V�,���z�}��s2�>��=�E�@��z�[�:D1�ں?G�j�*]�ꦦ̏%(���R�l���\E�$��}��oḟt?%H����>	�_d2۟��L��0!q��ٸ��ܷC�t�p)W)�9 \2?P����q+�l�RM���̈7	��y
�8w�j�hI��T�d]X��M���k��Ϳ�\R ��m�/��3�:���~ɉ�4se�0o��s�Ҥو$ST�a��ZD�ʤ
�;!�!L�Xޣی>5�e	dٻ-M���0&�HRԔ�+oR|:���s�z
ْt�ɏ�����)2VDi�B�r���x��~z-�l�g0ξ~9%�8�%FJE�.�(��Oڽ��آ�k�B*׀hB��σ4��C���%~q|~FAP����H�j7O�0ދ��{\3��%�cft˽&�$0����A�l��[f�-�������0���
��bB�! �:+�;���z�^P�ʶ��E6#���"����Vu����E��yV1Q�{)���\>��A��Nt�����̌�+zF�Az16G�Q��_*�V�U`���uȨ1�F��+^h���&��͌ �f<�h���Q����T �p|�B�Qw��T��!M�Ta;��*��-%Z0�9tWL#�D��޾L�2�8��ΰ�ܽ�y;4��֦���3�\��EY^pm�����H��+Kh��w�Zy |�>/P�Sבּ�(��eU�-�⧓I��bg�~;���C�z8
FlE6��t�WD7��ᙵ�c�99rݨNf�N{����GȉD����7"�R����>OoEq�Ԏ�P������]ƻ2���a_���"��v�1*w� %�ͯ���C)��Rp�ҝ4�XP�"������cQG�J}�G;d�x���\�P�i��������gbw��$0,:n�G!pA�����z&�xiOh�*��y�:���ie��6Y����x�B��ew��&��f �?0�C����*���$�k���s�w� ����]�JS|�
�y�v�.=��=�)�~��v)�ӯ����H���m�΁1�)�̒���Nb+����b~��ҒH�p��Z}s߈�FvInd� sp"x�2Wofo��Ռp]�k21��٣p�����ۤы��~ə���H �"��7�+���x��j]�1��=b��_-� q�G��+�qV���z��SJr����ˇ��(���YLO��^O9����Gă]�u��xfH.w�|���F�Pf�@��P�R����ax}�v��#������9�v�
 �{���n�$����h� "'��C~��gk�us�?���EB���R;��~I+Y3a�r_<��&��'�Ȗ�O�ܑ��mD��Ϣ:����ho��RnPJ���i_���:�ӿ�<BG��7$�\ŗi:!!�%r_��M�T$��\'Lx����m�hᴌ�Qn�$�h6H�4��;�����Q|������UE��[�Įq�sj���� �	;�Eq��4z���P@�#��3�r���坳�-}q�DN�o�e⬰���?�Q�����Ҝ:��/#��P�8��_�@��"!>�<N���G�W����NK��˱�!6�:�j�*;,\'���AH��j���/:H5��O>SU.'�d�=/��g�i�󌡦�NUEʉ�����dY'l����l�;� {�4�������@d��>�
�$bZ�D��-MI�7�J����7�xK��1�I�@u�ܗ��١��I�e{�斴j7ˡ�� �`Hl�
�%.���f

����M�D_%�SuO��������V��ut��-B�iƨ�t�`|��X0e��R�����eȚ��w�MOU������&��V�X��6ɏ+WY��<xwC�N�|��Ż���{+\�Tіzrf����
�d��^�Z��R^�G��>��N*��x:�-��YGNFf�M �7�Q�G :ѽ&7/0W�,�2υ�Ų���4��N5+��>�>	�u��F�2�R��Y�	Z��m�j4�su����$a��� �&=�����iU#ސp�J��-;s�J���%<9B��)aiN��C(h�PS�����}&6���Y��0A�+9(>`�s}w>s��qhƈ��̩�ky��˻�Uh�x{H��n�v�+�JOf0)�M���xx�؎�Jv���dP#�w��D���o��Ɉ�T�ֺH5 t�S���n�P�ͥHF�!5v�~@V7_G��5���K��_����&�~��]*�iG;&"oP�S9����/�G���.��	� Y�'n�%|�O͞��g{; ��+�g�,�$*�sOk��h�5ܴ.��ӡ�;��]i��\{L�[�"�ހ��"^������ו&�_>mw�uܶ\�u<��%�?�t��w혎6�ry�Z��!Οo�b�woj�P���3OZ9����k^��ӀT� ګ����M;�{�W���G9���8�1C��:�5@�e���}���v���ΟR?��9�#��/�e�ȫx���+ �O�������6�h ���!�]'ye��i��,�'*�,J����9�~>+b�r~ j����U=p͸K��t�ƽ�[©���-��v��/�bf3�p5sJ*)�f���plƖ`�D� �Z:cVo*=�/ϩ�3ȳ�������aB�E��%�����+���4u��>�lh{?�Kq�s��p*��IP0M���I�kC ����Mϡx�X-b��Ӕn6�,�"��h�����p<��k�CsXX��<j��)k�/b'⼍�v��-??�>I.��Ҕ�R���M�^ɑ#�|^3�f�>��[4f��L��Q��> {�-�Q	�?��m�h�����$��~R�>[��pU�츮����b��#��n��ҭ�Diyޘ��.���ȯ��sV�Ŷ\��v����<۔gC�����������?0�S4���>m��YB�v7��n�PQL �1��j*�8�FXq��JFi~y�)9���:b��9��ɀ��9����̦S��wX��t�j��fR1du�	�r~н��\��������Qƻ�Y���[��>��	7�����I��� ��=s�x�=ŭ�?ܺp[]-S���7�]��Il��&!Y�ğ^�b]^�:��6+�&﨓�j}X���,���z�9��q<]�"�pH�M^WT��6���sê?���C>P�x���@	����Mef$wS���V� �~塌�;�`:y]�6_$�zb�9I�8�`����%��� ����V-7��KQJ��]+���8���֧��n�E��H���ʰH�NdQ�i��`#���z��|������0�IC��0�v]�#��ڇߍn�~pf��U�2As-�?О�Tq.TGf����ВX�>b�?s������'l͢��o O������*�B�i�o����D�p66��)�e�j0��
r��7v˰>�?�Ͳ�?2�65�w�X��|tg[�ֺ��"N���D���3��m��&����vSY�*~�q�����Y!_��d����d�)M(�J��p�S��%p��XI��;��p��^��Q9�`*���%���P�+R������B|�V��'jkl[���h�� �%dx\z�;�F0̽q-��Hy���?��Kk���?�Aa���(��>�M��G�H���h�;~X�y#A0���+��-�!.Y7>���e�����Z�`\��Na}��FWw1[c�07���=o:��	h�c�w�yl�9��X�Ћc�iщi����"�6�O7wJ��XG���t��\<`ۺ�+n��U��L�#��҈�>�T�"w<M�Ba8�h��2�A�a�_o�7�����j�dD�<;m��B�[�B��a��\|�ƍs`�i�p+����:Jk�TB��CAO&�r4��:7g?vYI��M�G[���۱�Z4}B"��Ϫ�e�'��.Ɖ����Ika �x�[�=F���,f�,}7��v�n3�=�{zv$�F��}��I��v�e�c�b�!7o�*�֌.�K���\t �Fl��U��2y{M��. U4_��z�0+�q&*�L�Ux�XX&�ﮨ]�-��[����/�
�d��)B�L4od�_I��Hur����_� ?�1|�8x� 0w=kLlv�R8H�V��q��=/QU%����b-`
�/g+���u�ܦ�n:�(]�aP�x#�(`촐�X�QP`�7LRa)���iM3.�"�&?]	z
k=|=��(&9-�j{#�N�f��m%���!ESZ��Rl�Xq�P����C�F4s�65�1Cɨ�H�����f֛���׎�3n�gHq�/�}����꿕�?�-���)�ͻ��ms�6�:3,l"�1-�
Sԓ�'��eWK���CI����h��.�+Ò�=x�G�>ʲ�r�M�:���;�Ƀ3�������d*$E��7���+ ~.
�!и_��Mi��y��w�������V�}�qy�k�#I2���}nU,f���Ֆ/��a`�7�M�}�+pJ;P�������m��b�	�b�`��Gh��/��g�C�.�]������Z�<��B�s��ʤ�˸��y�
����]F��E2�08zc���b�"	9������_���U�����h�`����.��HeTC�m�����N�=��r0��g�݃�jʕ���h��Ěj��y��Ka��n\�s�E+��c��,A������Q>��;�1^.-߽}��W�+XOH-�:�A�-W��a���tþ,�F��WF\�mY�Ko�SG�IYbul��i� :��D����]��U<�5��3,���'����lL|���C|��*�S�^��0�[-��[ER���9�N�#�)`R5-��?�X�o����>;ʉ�`f�/y`�'Je��EPh�\4e�E�S�zإ���Z]@1�ѥç�͈ڰx�Dz�Of� ��܈d���P1$M�[?���*Q�
�����֋�0t���CU	; 	ǀDS�&K���&8��NY�m�F�6d��"lZ��M�m,��B�R+����#���c��J�"��OT�ڇ2]#�O����`.��_�H��2]3���|�g�q�Ȣ���3|���^��nL�Lh;�h����l4T���2�\���;N�1��4 ����S��Td�j˽�ƙD+A aL��@&-������Nţ3�v�H[R7k�"��"2!,\��f5�qϬ��^#��u��*6s�Qs��P�1_�I�T�6���V�ce��,��J��0�܎�bG�KG�3"��7���h�Z�.{q�Yן��T*��e��9�~q�%�����ے���??ܪ �;q۴����I�iȒ�������� dM�:�'�Ľ��kk[��ւ��$ĄG�$>�?����h((~p�A��RTi� p\&ox�E3�k�����4�K�=X1%��������20��TS=�F����&�$Y�7F��g��A,�#\�fǲO�=X���ET�0�P�k�{'߭��pg~�a����F����3�Y&i��T\.�Cf�ŵ�o��r7'��H���5?yb�ǁ��p����f������>�S���P}xU�*F���y&���$�]o����wgx d%���/ϡ��i�I,�]��b}G�p1/'�Cy�c��iA�h<�ɽJ|�d�Ԫ�Ii]_}z�4="W���(����:�����m�����^��x�Wl�b����蹟�����q��� ��\�)��w3����%T�H�e7�gP!嶟�peu��b��0��p�dԀ��<�1[��e( Tdo��w��"0����{L�|_��$�d �B��Q��1�$��=��ت�/�\�͕y��Jͽ�1%)�&�c���=>:bd �Kv�(t!,�e~Y�qe�3N�*_>/|/W﵄�4K�w����K�g�--��E��_�����\-S1陕;k'x�$���4z����X�*���I^0�:%�3�[j�$�H!��Z��cB��.2j���~.}�Z?E���h���ae��غ]�\��UE��T��^o�4�b@X��!�ix2�B�.]��%5�2��"(�_�j�v��iy����R�<�>ѳ�L��Ɯ�)�y�	\�{�aD�APD?L�Ԏo���m������r:�R���!�\y��X�W�hD� �!�oql��j��.�@�RL���^O�F�q�&��g�P#��uq�Xa�f~��*Cȁ(;;@��4�3lR|(��tM1L6���:�����*�5~*+�J���!��a�9D�%	�
�=-��Pg��߼����O'6̏o��)۴��X��+NP �w�G|	<�Vߣm�dr~��/�n�wn&b,�(�g_|s�8�㈁��0���\�U�bxkw��:��H�iP�5m=u�טy�Vi�4�ì��e��&҂�:7��^%�,h���=���y�>���L#��o�P+������zq�V��?��yޱ�݃8��>
�q�^��*��R��6D����zy��a�YJ�8�wh��f%��1::KҾ�	V�.[�[��Io�6��}�:K���՜=����2o�~�l�0�E�'��G�"a�e��鵞�S���?���nqt�5~���,JdOa*���A-�n��3����|1�G�W5qے��h��o��0���Y��B�N�C�B�٨Kn��1�y���BU��ָO��>��t�_S���!eo�Ϳ�x$�?��]`�&���{�}�
�~;�H����}j�3�[9�t���93�a邚�}�����	[7#"�)��4���ll��L3��b^&fb�s����GBx*�_��K�*	B��Kf1)�Sɖf�H�K��ݝ�I�?s����k
?��yr׌��O��[8�w9��7�6} ��~ �Vf��)'�������tZ�XB95n�K�c�4J�يMI�B�nb1�&�b�BG�1Sx�l��xI��a��D]Ԩ<V+CXh] f��4�����|{,.��&�{c,���&ȁt�}��$��}�9�c�Y�j�iuR��Yׅ�I��M�z�bm��ЈWA&�t�&���t�O��a�(����^)��h�uW{��$��ہ�,%�Ɗa8ȿ�6�-{fۈ�܈��fTu�vvt�o wϓθ�{]�M���Q}�N��}��`럷#��,��$����&3��{0x#�/r�F��ѿs����u��ql�?j���o���[������J��%��Ө�d%Gn��x��/��\g��n	�OL��������DT��e��s.������Ee;�z�e��D��g A�gdz��X���-����Bix�$��>����^���{ʫ���"*�	����҄�I���]�h�ɺ�z��/�Y!��SbwY��]�����',���߄�+1<֡S�V�U�����YR=u���@5w�mdS~�����bA���AH�E����� p�Zq�V�,2�ꉫy�7���8���rì�yj{�4ٝL���%
qs�z0Vq8��#(�#��j,F��v��Om+̝B�P�z���\\�^�L��N!�[ZzJqU��j�j�fh��(G �ِ����+8Xd��Cܝ�c��\)������:�N�Z'��Z�p�S����Z�M��1��R$��N��ߦ��ī�%ʺ!�\(u��I)6��q�~�S��q�K�����<�(�4�A�s�E�I�T�v�]^U5���bŏ5]8X��R};��+� zX�6�.�7��Q���f�;�	a��F�a�h��,���y@~Hf�����X����M��8[�U���۲Qc>*�}�BlB4�#���g�Cr��=sq�����Uҧ�p��Y7�d�tڪ1��L������
Q?t!��r��E`��ak�{t����T@��'m�u�hPݭd���(&��RO]Yg�4J�g@�i3a�j͹���B��:=T,3��NX5 �i	5�*�!U�r�ǣ�AއUG�����������T�Pٗ���d��Gղ�`	����^(��)[*R��q[t2 � ��U������@7$f��ޣ��iĴ^<�-�UN�����r����R�~����|1a�D|(p�Z�dj���������o���l@���лgr��#�
�{��9�d5ļՑ��s�M��܇��ƴ(=u���QKl[�^�>�!h��L���Xq8��n��lP��	������?��>YT,!;o��O����CU���|�ql�t��c2�h���c<�� f��7�˶�s���ѷ\��n��M�Bwbl���Q^k��q�f�䍃n�?uH�"��\�0�>FbhTM\�p]�;���&O�l/��G3�ad�+f\OO�
7�Xq���e���-��ۙ�Y*�(υ�Z�Iyx��{U�b&6�4[�x�M��aĲ���y��M�"A2FN�����𐂷P(e}Y���:�*�Ƣ���whZ9a5TO���x,B-��~����оM
�����.�F�6�L��fp�$�ShWq���,��ن�����'�g� N���-G������h+�8�����m��%�$�[���.�����8{ʀ���&-y��&�#*�H��	�@������f��7O�pgO�|,�ƽ,����Z��=�e��X�|K�@$����Uv�֦墛�QG�� 6����k�J^c��4h-h�R��� �@ �:��z� �]e��w���D�Ks�>��-�\�7�yc����>�aq���/�ð��r[r�	�A��f^�E�k�|�7(�:��U�-�kr�:��F��9Uւ�1kB�l���4ұ�s�y���~kw�Q��`�GP���g�����Z�����ض7����� �T�PF��B�>��M�͋�.I�A�N.K�dī�Y��Hp���.��9@�Ϡ��'�7`�Jۛ�77��Ût�`���s�7���ȟI��U:�g�+�1Nq�B ]���M�RdF	�+��hTC�0����j�������l a�|��n`�E�>[ٞΡL9��̌���}d>�
i�%��P{R\n�]�K���jr]�ep�=d�d{�۴0⸥QD���w��u7�0����?�I&�pfԜ����b����R�����8�	����?b�ޤ�]{XWѐdj�'sl}�sQf�?�(�*����P����"F�) �&5_�R�s"-�oGa��;�BhN�K�#D��So������]�I���2��Z�+�py�n@z?J(�!��~뱚�U�s��mD+��KM�%����͂�,$��i�㣟��kK��mµ�}���=����(��C�0X&8�|%P�/�bH^=L~I�l��5�hD�z��������|(�a��WH^��޴�H��H�x	��lۀ�����x��EN���Xr�>���;��2������\�q���̎u�u^T�8��~�=Dg�	�ǥ�$�?�1C�d:n$$����MŸ�|F�����0 �)�1��8w��7�ګY�+xL����V��,2ķ�@���1M�_��4��(S�r����}���O�"�tX��e�P��9G��zf��dX�N*����~�1�B�O�N��H����j{l���.d�Ц�����3���NZأ�~�������j���~��I����I|w6���>���N�asJĩw���N���#,\��QN�k5�����s�#��8��3��V·�����j#�,`R�*�,�Gb�;=�Z�ǀL�D�;,#�q@�]SVCJ��>Xj�}J�=�C/<�04/I�����ИQ���H�N���]���x��B����c/Й#=!F��Wg��ͪ���,����Ώͣz��c�	*]��]����'e�p3p��ȅ\,�L7�fQᦢ�E��rꊺ��lI׍q�-��֎�}��n���|�^~Cr넜M�$#��M�dJz�d���rܙet�Vs���s�G��}\�����x(��O��*[:D}0$���\Bf�& l�I�xչ�vm(H����x��(����m�{���lJE����C�u7`��Z*��Y�Xn3��0�N�jPK����s!��V kB��{:��!+�`�e�v�0է��\{������߾��o�5�Tg '�h�?͒]��E.����-Q�3м��%���>������2�w�Co�k)j@��)
}_yoLL�9#]�����*�����45�*�IKi's�[B§S��=�\1�,��ܩ�h�H��B�<V������{�6-�7+jt\�2�;_���K�3�G�Lelϣ�e׊O(p��^�������fN�/�y��dX_=��g�7k��] �a���=^i��!B�	���O鉃�@闓�:N�-S+�S?�{9Q/�`/��=��{z�ԨX�4JT�������%ޖٯ���nD�w�'���}��뉻]K�@����>��1�38)Ť˿���s|�HѦJg<C�K��;�v(Kz,����D`�ݤ�8Q�~��싕2>�n����V�FqÁs�E%9��K�α�}�4Ƀ�X!� ^�(���77=���ɩ"�Hc�C�rK"���?	����,��K�a�|��8/�������:_��W*������0��P)+����8V�d��<��iJ���\�2��7��IVS��f$^�!�>9�;�Ƒsm�#�H�M�_;�0�@�Y,��G���ĸu,lW�GL�j���zψ�&Z�KB����駰
�}�lˠ��~]�����̬O3b��e�5�}��<�ӕP�����FN��ʤ��jO�;m�2�Έ��aX�*c��O��J������gK���r��+�K�wGh[?{�D{��	�wQ��4���r�g0_V����R�C���0��0��SŔ�n�X�/��ۨ�e�}��n&D�x�������s�X*����B<��+�[��G��E��k��}���i�Ohqo��Ԓ���1Աz�-��泃9p��bQ��6)OO�%(*k���} ��SE�t�l��:S,Z
�?�7�F'��A�����{O=FɅH쉓��2�}��*O�$ ܺnT/���')�Af�:�F���F���ȫ���.�����aO���3�#$�U�z�e�#�N�ob�zxm_��O�%��as3�{�Zt���m!(vT�L9g"�LO��-�d�
K��&�o�� ,r?�m�K�¸
i[�\��ke;Y�m{n;HC>]+��������W5���Z+���6��/���*h�-w���?��2�ߘI�����piĄCx3���vڑ$Vf6�������+�Q�w3^ ���cwE�OX�R�� UJ-��� 7�����2�g��l�>�YUڎ�wnP@7[�[�e%�	��ٵp��Aϸ���Ijʄ�J'������h�z|N�&�/�G��4s[���I����c��+��M<��/!��)hp�~\���B?t���·Ķ�z<�tW �u9���:�:9[xf����,sbfC�dWޫm�äL�VgL��IO:��[�$������l5��[��6���o�ƶcP��[[8Ι���6Y��.���ǟ_�$�룇���/� ���떼��n̺=�-#���������4����'�8�|.u=�{2z,g�%V�e@�h"�4��PRp��2�b�N~�6�T9�����s7�|��Mע��a�DO}�u�!��	îc��j�������{�����&�)�k���̷�T��#R����	?�gD�EB�I�S�/�"M8���uڏ�r���ɟ�x$�z��Kz!�9�[X}r
��C! �͒d�9/�(bzF��V�e�/) _��Se*Swzi;g%�v�ƶ*��l�nN-�f�0�	�&Ef4�L�.�)f56M7�"���iȉ;d�%6��0��y�L��~06��{�E;�R���tb�`�7�F�1�RTS����#8D�`Z?.���ǩ�8�ҡp�D�f�H��4���Z���s�K�!��� ^:�e3��&"��)x�1×q�i��eVG"�SX��l[�#���c
q�]5��'J�Q�C��A0�	b]
B8�zr�L5P1�j
�;��͈�Qh�����}���%8�K}�o�JM�%y,u���	u��T�OQ��EE|uSa#��D��S�}3 ���v"Y�A婯\\� ��� �|#��M�yB�a<��kt�k���e�߹2��L0���e�N�LSw[4��h��q�Eo��+������s��[�9�s�����&�4,X�oZ��{)/�y��xL�ZS���V@.O�њA���ȵ),X����=1ꢆP��>�sQ���w��p3�O���Mn#dy�)K���3�$Tz����\��ǋՕ҈Cn��a��^����]��V<A0�&������vC�� ל�׏���>R�)s�,�Sߝݩ����ETu���#���8�F $��v�aj��S���St��:���9���0��m�1��oW33bo���|�^�la�<��@��.ˋ����V'o�KHo��6| �����|^�N���E����U�T����X�\� Y��K��fJF딆@R��D+�nnXr��'D��("ǖ�v�|�w��kl�ض��;��Oq�_�_�����]� �;�7g9���r�C����]/�7�{�a�&�<ƈ���_���s�9�L7Z����r!$�NTL��*�#9�c5D-��u:KW;i���w����j4��r$]�1hve���������rv��p1�ú^Z_f�*��o�I<�~K
Z��� ����G�Xt�����P�5�Pf�iUi[��f�H��#SŬ���	�[X:4��L����~����fY�/޿>p_P��k��I� �$�M���nz��Y�
@k}�����h��ۥm�ƣ��Ax�o����#��94��q3�ܝ���R�P�b��3��`��G^r���#, �>�� ���܎��&Xߩ�uE~����| ~�/P�5j��Z�Y&����]1�"~��P�M��S��8%�g����nj֥��#�񇽺����r����jҨ~6��H��s�xцȒP�0�b.�����Q�S��#�F`صX+w^w1��Go�z�@L�-}9���oe���h[��,Q,� �/S�^.<�P��T�x��������0��N�3�Fu!����*�&(Z1�0�R������X���E
o�??�����m�G���2����b��V(<������vs�~�,��SI'1v��-��z�=�gT&����c��+G�j�|��Dp<�G�7���Cʦ:1��N��d�~[����'�=*n�/S�d�����,�<�8`y��%-�w��A� V��ݹ<�T��W���J�*y����م�Zb�������N�@��[������n�9Q�/��f����כ�P<��)��2��$�Ԇ��Pw�-���Z�v�������r���9@ۻq�0u�����A�������^w���G�A��{d3���@`k��7���O�p�è��o��.1�����z��1�S7=�>�^ ��4��SB"�t�I/M%�T"d���b7$�,{�&�̟#�5��o��R����~9��յ�XEg��0`8��hj��hU�}/�7Mt����82��T���&������J�P��_�[�J��вذT�����R�A����6zkC��c�i�Q`j�,�Te\GR��"��)���Y ����]<���eJ^م��c>nc=w>V|���odO7 � J+DT�;�����b:�&,\���/�����������A�o��r����GrA�w��؃��8@.s�C�t/ç|����/��#D�U�6q�;�L���i-���!Y�0�x�~5O_C>K��Y�(��� ԡRoe{���9��|��&VW��O�m�'������E��N�S�߮��&��Y��3W�nZ�ƒk}������g庪�'�47�0�}q6<�~��j�!|�W�g/[��1hFB(�����IF�'xQr��èC�Ym�Wn��¬P�W�")qT�TM}:s�f�u.b� �'���(�Q���)�m��#"���?��m���{b�"����=qn�PX���éQ7�vh�yֿO��&�hЃѐ�&��U�TQ�_�e�cCf��I�B-��fў i'����N�*׳��܉����L��K�Gp�UI�t���*� +���-�/��M�\$@�Vv.ף��Ƽ����s���T��4�>TM)/��K���R���(�U��<��M��g�{���}ׁ���Vi���^��s=�j���u�E�s����T�cgȴ]�[aEo"��)Q������і��4�83~=?S!�e��uZ��j�ë��P�ʲA@�`]�h:DP�EG�U�����
��r��[��:K�Ԋ���غᬪ�F�����z��a	B�H�4�+9'�jw��=�	l\�.�%%��[�`��q_2��5ʩ �K�f��M�O(aW;���נ�ļ�$���Y\F��h�F4��}������|�u�hxw<��HfW�(��	�0`���Y/.�5��_fmk�	_�0����9�7�wk������v2��5a��_19��0�E0^K�j}I�u�#y���3U�����N7��j�t���K�jM�@�p�QC�F	��PKO�g��ƓD9�N��3 �H7�,���@�̏^	|��9{��eP�{1Fqs�����W��W��F��(���Nf���;����|�&�������zڟ�v�B��?�&JT� ]����}PJ������u`Ueh�N���Ԡ5�ZLlu<8��� ?]�ht��n��Lj�+��T�
&�@�Ym�t3�����;K�$FT��b8J���x�H_���1-��q �K��8��::C3}��:mj�SuӖ^G���ր"�|F���YoF���ͱ>�(�5�7O���R1��+�\�ѧ�ɪ��.���a�D���W��+zœ��(�/� e��I��O�̤��+�JT��<≄?C|���0i,�=�OL,��=�[6��Gq�v��a�>�W>�It�:[MYu�~w�*A[��l��<���0W!LT.��6�۾e��-���a0���VۭN&�2 d�Bc�ϑB_�,�z1���g=}�i�;Ax�"�k>6�>��L���}ngp�K��w9%����4L��)%a�@�z����sb�2)k�%Y��f��?7,Cۯ�2P�A�I�W]S��F�$����/��4��H1{��LH�ja�)Q�%��-ʍ/Ń���FF?U���Ǻcp��1|w�z_�AqE�5�+�@�s�]�E�
��\r̓vF�Φ�e��H��?B�����j�,���L3F{��dD�x�!!���Hյk$*��#��̕b�[-%#�|����3��\Xp����K�V�'j?��싑�?n��m>��O'�DpC��Z�����Q�f����z��?����%	E+����箨;~�컜�؎�O��s��7L��lGsM.�6�q 	�Cv %v��;�Ι��ٶ�A|��A&��Q2{'ɾ������~�!�+~��7O~�6Z�G���j�W�%1��"<���<��t���=oL<�L�Dw>`�����>ΜN'>R�ҙ��4]5�rU���*48�(�t���(�F���ȇ	�!���2� �6sN���i�蝽���ѝ�Q�ņ�K1��ߛ��+DP���q���E:p�����H���',�A�����Ė/�7��c��;�^%���c`be"b�5v-�{a׋�A���H��Q[�7�N�]QC�c��@���ݓ�L/�����a�U���f�mq�����R�"���1(���hW
g�_=�@�&���]�}@�v��+���Ujp|�侇�O��~�V$�L��$b	��&m��#B^yؚ���w��x�\��R�����K�5V�A_%����"�g�Xi�k8�^�x�b(�K� pV���h+Ux�_uS!��ݫz2~Q��_v�N �g���Q��L�๕���e�4E���u�~�[�iVx�R���V�Λ��S���m&j ��=�+Em����G� X{�?Go�9��h䡱�y.qq�"ـi��߈~"���o�Q	����f�D=lE��h�1�ba� *�ۋ���W��	����oL�8&��Ng�yRڍX��O��ZU��9�͆�g���s��,��������Nobx�p����T��<*r��,����"K��Z��n�C8�x�r�`����Bt7��	LS0�2�۟|<ȵL79���&���~�|�XI98���4W�?ú���~C�=O����d�����hPW
��`�!D�9aL�X��H�����mZرZ���g�����:�ɗd��-�H6Q�ƻ���sۻ`El�M�s�v�W�;�d;5���>2l
��DV�$�L�ԓk�k�ۧ�`��#�����0F��(;�{U��y:23��] A�W�&�_ϝ1����<\�ɩ��r��U��x��f-���b�/ g��!|���xY�q��Ԯ���^Y�pu��4p����-8�`�r�J�� *#L��ҿ$D8s� p���&�}4+�{#߆5�5x{��ag9f�~yҌg8HE[ⴻ����F� q��"p��e�[��^��D�W,��*�.�Ut=�2"L5ޡз��b2�#�n��;7Rmkx\s<��vq�P� �����������σg�h/��J��l�!��烙^�E����6]�'C+_x�h�:ȶ��^��ƍB��/�i�N�¼�e�[�K[1���=���F ��7L��sZ�N�_q�;����\�b���B%���,�~e��ӕ�f�α��Z�o������Y��"�`�pU`w�P���rX����E	�&���SO
ݍ�L��~ZQiQ�[�W�E�H�g�0St�p�V�H�H�S�0&$篴��1�Տ�G�Zs��:*]����ǹF�0��:���U�eA�r�����E�S�f�XE�������+�U�^��=Z�Oڛ����	��D�˲3@a24�~�Ss�/J���D��t'������Ե��hW�?	����6W9���H�Z��VJN�.@+��!���3�/�9&�����*��H]���E�H���zQEeK��I%�Cy�@���.娰�sY�n�K���|��Cp*��O����Qj��L���ԍ�t�l���f��9U���SߩǣԒs��}�'ԉE�8ӓ�!�uH�@ĲPP}u�2GU��O��}٩�Ph�Y	!?}�H��>A���|Y)��<�I�hj|���W&ַ�r<���;�5�\�
��`꯵6�v=�?Y	�mw0�y-$#�t훩�	x��x��s+�ß�{���ݤH���NVW��z峊P�5��m�����R�!{�R�[��?�jx�PcΑ���k:?����!ăܮ�鰜m>@<m��� ���Vr��H���o�,��%�6��P��S��E���}4�;�u��= �U��j"�A�CQ��;�8��Ԡ�*��[��o\��z��ٕH�*>�!�}ɦC�Li;ڗ��� �G�a�h�>q��M�����;�2M�͔�l(�ۮ
'D�C��u��2���ՙ3{�I�Φ��%l۠����G��]t#d5K�����#���.���غH�ᱽ{�
�b�� �F�p���x����ۛ/���7�6a 0ؔ#�^��d�bpi��^��L�_��ЫRN6��ܰlr6�/��Uk2�Owъ�=<�l�L�c��^�s��/�;�=F<�b�.�)~��S�opS����l�c�E���%o0)m�*�i�R%�i�qT|��t(�Bpu��,M	�����L��&�TE"D�K��iV���*|�aN���V�v.�/	�JHx�|#I\�LV��h�Ex�������D���:����ю_P�F�֨%)�����H��Y"cP��Mf�v��0��� Q`������8q�ʸ�����2�y�`��bfm�ͦ蘗@»��� �<��|/ݟ��R ���U/=�۵Dj�Dd��X���L~�ޗ���c���ˍ�q���&�ԑ���D���2��Y��=�nPL���ቝ-�֪6ٯ��i~���?��f�?�j\����8��:/x��ʉ�r��ůq���a��(�G�|������qz����Ƭ�X�$���J�r<s�d��!�gE� [��"ֻ��C���6)8�:��'<-z��C����ՄS,z�υ���R�gЖ�=4�`G'v� _[��{Л2f��q�_�̎R$(
����qz�Z�k�)��Ð�k�|�C����4���=��45���fHV�� (J~v�GfH��dl���59	 B�	�I�p�R�{��lM�K�g{O�LN�\�p���L�L�*P7�T�e��5��'�����e�2���2�d�J��$�˲��[N�K�w��L�gz��8$�ns�2}s]���ii����)��Ne֠�nص}o^�ͱ��,ꔢ�]W߼����,����T������gMdc�tn�uF�'2���oE��?����䫓����*����*��?4�;���#�G�K�V�w�����T���%�zyr���<�=
B{�!�_�@P��|���i��V��b�FRh�����,�/EF`��O�����vp�����'-y�S��ڻc�y��[�VhP���CVW�MH+�W��k����v�u���I�<��֋͘�a&=�lHh��`�p�/@G$�Y�x��Q�&��c(��V��
C�6@�7�T���h���|r�,�?R�!��7��L
�K���-�6�� ���4b�}�ڥ�D�J�6;nTi��~����:��}�

��PEU���\ΰ�uv��@m9)f���oW� "�	�@��h!0�%A��O�â:�(�<�6$������� ��Y�O�k�ԇ��c��$ғ�|v����9�[�F�m�[��n�{b)�ry��vR��ND���w8��UP0�/M����}#�[d	�Q�����q�����F�(������/��a��Ghr�ԗ�9�HA�����DfC�r��󓙨��:D�c��k0q>��fI��+�=K�y ^����ƞo)��<'Ǜ�	f~z�:�׽�o��u��dE�`���ْ����(=<'oBI�������?!��tD����6�}rzk���ϋ�@<u���ȇ��ҷ�}"�T�XJa�.����{.�����O���I��
4�X[\(Cqk�~Xy�����Z�G�{��+�VP9�u���gC�tz�N:�Ո
<gIT�;1�!�����g�ID� �.5��	9T�#��n#KB�ynL���RZKB�<�Wc>L�*@.��z0"^>�D���NH1� ��SW���("��z�&���S���ݖ�v�J�)O��փ#�1�Yq�1�W���#D���پ�7H�FV��gw�Az���]w�l���r֯(8aX��$�fʁ�g9�tb���Mӑ |~>�j�qJ�@`��{�K��ͫ�H�$�%�Cl��&#}7:��9uNXj)�)�5w��Y�{CT,\+x�+"�G�$����\]����Kz�
u� ���c/Y����?�l�#r�R��̨�n,�&)��]�Z ��i�Jڅcd.6���p�4�5��U�Ȁ�
�d��~?Xrͽý�C������/� ����x��8��Հ��;6}<�mח���>D!u�P=e�(*���"5c~+Rb�����#}�a��lR���=&��g��5�EG(�8�IV��f=[����qg)?�f��u�1�y���;&f/V��wD��8�JKM5��*���)V�c7�=�<؊�^��ҧ�ch�b�
���V��n�{�W�l��9�zE<<!�
5c�
�
���o��0x���*�E?�
ڷʫ�!Ӈ����/��L�4J�jȴ�����X_�YJ�|����1wO��]��k���P�?��~�50�% ���'�����办��ٖ�s�K�Y�j��q����gd�&�f_vV>���q��k�{m��_}�z�}�h��ŷ�h��}gGC�N��ѩ���Q��@�y3Z�?��n�B�Sw��B����Pw�o�I���&$���L���瞱�3î$K!s���8��mݝ��l	��^PP��@�3Z����6;bL�J�PB=F�A���<�tg��5C	�rq���3�п��]�eq��p�8}\�%W���3F oA�S�W���R�<��.2v��X�j?��5�\��Yq�m̋'���<�^03%4����=۞���(C��%S�iP���O}4�<3/oc�I����QsV�3$�i7�V���^(����>k (T��V��׊�H�����l�~��ش3�2Cһ"�躂����
�=u]�~�R^��-���	�u_�`���p�?4#x� u�5�2m�[�+'���d훧-��LD���>��cz{�:�v�k�Հ�_ջF}�S�������%w<�i;;�n��7r���B�	:�������Fۤr����"�^��݅�����@~�L�6�ɚ)�Q���#��������䭱\:�Y��-'�vFJ����r�=�Ut�Q�d��&�u�.15�9)�[�,��4P�̩~�& 1F�y���Y"B;��]BA�m��K?ј
E���N��M跮�Ⳛ֛26�����ry?�>����� �䈉|�k���B�:"6+��z���ex������)\�y�O@)��Md�;�x�PO|>�Z��T�{���XI����P}Z�V��h����8˃���O���ߏ����¬��#7}�� 6�1i�-�$�W 54�9��7�FZ\�&�`�I.���'����"������7��MPr¬SC���b�j�r>��#P<F��r�;�8����/�G�%�,��գ0Vf�E5�FhF�N�3W�����q���%���m=6�u\ޜZ�6sFN��~i��2�4����waH-6t<]��D�sbi̺̝\YT�7�����V^��A_���%�0F�s���F��~���r���_�*�\�4"Y�}6��{Po�=
�n����Ǥ�_1_�NC��'^ ���d%�l��9�1w��z��y���g�5��p&�?Q�Ö�[�A��9U�h����G�y��V��Rgy���0b 8�Mg���_���
W&�.%{���(-���궹<\�F��"�:��vTBطƄܴsmV��Sh����!����_��e3���>�!vNX���G�ҫg�%�]�u�Ż���EGwUñ��F\Y5��P����t6����%p���'����&�؝M�`�`�k�f~���#k#/ �o�DW(�&�.�L��{�1��w�\��@��:�Tg�~�:t'�O���+β/y����.h�:�DHL}1Ff��:���v)��8UH���3�_�^k_E�6Rʀ��0��������0F��I{�ڭ%���OeQ��E��^�l��D�ʀ�L�04l5Ă�b�p��p=��rnb<���5��>x�.��y�l�=PZ��R��[2�<��㮻b�,j����o�|o�#�`谉���,<�B9|�`��(3�{RQq���KTj\Lv]�#��l�9\�Sg�p�bX�����5����4�(8����V�ۇ��Q�}�鐏�>��_R����
��~FD�9{�43���.cPv��+i�.����FG�%�KS���ҹ�\%�`�ꮗf;����\�7o������_t����C��H!�I��]I�Siq
*\p�P���D|����Dx����nV�N��F�}t1�7%,���:���+
-�%�g��ӤbGy����1`j���@<kP3G;�[w��/��rh�p�e>Jy" ;`�M���Ñ�������B�����`����=����Zŉee�v��*�P(��tLA*u;�����}8�/��C�.vW�_��	�nSҡ�0�����ʗ� ,�aw<q�vջe\�o
ϲ(�]�7B��Ҡ[f���ؚ�8��qJ{1ح���w%/��8�aP�{BU���]�M;�M!��YoS��Xķ6�CW�%���1�N�j`;��0��r/�w�`/�j�ן�<�d���/��4���W( ,�X��7��&Ѳ�Y�����ʨ_�^�dsN�����|i�� �,� `��B�ߪ��5S����s$L=-�Md�J�??�n ��2z����lm�% ������� �I:WC�z�=���d�y�A���?�{����N��α/��Af�XA��m5u�Əs�wMyv�뗌캮�aKV�̯0ٲ��������RMh���-C.l�QLJ T 0��A/b������f"�j�8�ꦪ�:�K�P�g��S�%k�;��嫖�~�Y��n����}c�OІ�h�)mZpSAX�)��|`����OSA�d�y}Xذ��z+�C��p~e98!��������1a�(�01��|j���)	�"#gt(��/s�y��M����k;�ܼ�k�_��=]������Ø� ������!+�H/�^_1��,l �S��"��`f�di�)���"ч�% 3��aG�4~?]j��������$�j��ķ���l&�n��%Wxd��b��g�I%��z��v/�呶H~�H�f_Hyx(�q�~;���`�N�E��r��x�S�z3jA�E��^`P�ʽ�J�	B�=�c}�m��v �8�Yk$�9 e:�\���қ�r�fRv����Z[i���e��L��:Ay����Щ�2<u�Y�
���ly�{=�[4�uۼ�ZxD���婬5s$[8��½�2��H�o_-@�����؇��Ď���k�
��gv+Y`�X���#eݡZ��uV��o�U���!�fC������5j4/�����u����U����m�H���Q�"֋~ކc���0�DܗJ}&n��8��f���*����s��Ӎ/û���V��s�C�"߲ ry鋰8���9ium�����x4��ҖM�t�C>O�[��̀�'����>��t4��҆���<��gL��h��'����^�X��̚OJH&3_��F����_ן�\��+�+y�`��G�|Y�b[�#=i��^�L��Ǣ��s;�ʁ#�m$߂,�2V��;��]�#�,E@���$�^���;��������3I�9d8.B��ߛ?*��}�Բ<�m ��m��ʽΤ� +�Ji/��mN�QX��{qb5�C!q���]]��M.���}��vcҙ6�p�3�}0:q�o���^o�c��ƭD ���k=��L�5�~ȣ�	����U|:4��k0��*�`����(���e�m�m�o�	��c���h����p�� �v��ꞲpkV���K�����$0_R�Q�'�R�B ���'�g�������� ���R+E�����),�`5�	MK���E���˯�P�g�u�I6~*UJ���-��<c ����K\4[jnb:=�!�:���-V3[��Z�!R;B����4����-ܣ��qH򠝑Ը�̊w�
�D0EW���`�2�hm �R(����q_
}��36E��S|�)�_�<��||�D�T-��6N�L�G����5DJz�$O5b⨃�Q�Y����G�c���C&��S��"DC�̬�����;ۂ3�fS�թR[�#���l�U.�%����1�e>|Ll�)ˤ���6���M' @
�vxS�MX��MA߻�7M���ۮSb��<��Җ��z�[��~9	g�����ai���1���D�_�T������}� am�	�ޔ����+�6���t��WQL���؉jBZ�^�(5����r��n��e���3˃�h��n������<�N����z���B��M�޽�0�PG|�,�EI��!vÉA$��q�y]�P0�9��o'�\��%)�M�����E��Q�l���D���Q��[��V4�YzX��,g���}��i�m��+�XZѧ��4׏w��H�B�03
�/�7;�۞�̇�`]�x�Wxޜu���E^�8�..1�eA�!*����u��6���*��r��;����s�|�2���"�sQ��J>1Qȑ�
��pa�D��WX�0�6�Ƴ���p�
���~>E'��˞�d5��ݓW7Mx�/C|�O(Х�8��=�^*�kIAtS��	/ʉ��@��S���9G��?��/�e�ݔr}�Ԉ�1'����&B�hh=�5sn����ع.̄��EWD{�Re�Ó�����)L���A(�堨3�����`�UU�Oir�ꛮ��ܿ{%���B2�$�[)�6Z!z�2k�s˷�Z�� ��~YU�e���{����){�>' �E �������L$�9}�;�VO�ss������Ynv|iO��a�㐮���N�[�Fʛ=�;�gt�?K4��ػj�i֋��#� �G�O�yd�Tw� ��5-�.�7?��;��(q�}��3��/�~�yp�8�O״�	l�呧S��A
�Ҟ�=SUpJ���^WB��QB	�>zEp���@p�Gj�k�Ս>uy�l������=DB.7��(�����<r�1|������mXn������z���DM����	RhQȉLn�>�5�i���?��3�:��1Eێh���AOo� ��9�K't�kS\J	֨�j����\n����=�I&�:�q�K�Q�_�)W;��z���3I{j!�����tax��@B��w�a �3����)��FNE��(�����\�N�;z�R0id�E'\�Ļ����ؤ�Y�:�<wbi�G�� 3��h�U����NR9��@���S������&^,��_�5;8Nn�!��l'~��C?��/��r��{S�0Vd�U��4_%�4
�:o��&�
�����_�?��#t��~�޴���R��Ts"��Wf�Lv�/�a7���֎!�^{�EmQ�w*q�`������hl&��l�E<<!�%�認?.N��-/HY
K�ZkB��@�d"X���oYӿj�3ڜ/̩麇z�6ʰXt1�Cƪ��s�s��Od5�.h��\�o�6Q�خ\C,lI��I�磋����W�m��1xu�\�`�����f�f�+�Q�q�����Y�ܞ�ZQ*����_��?�j�g�"��(�<�<Ϛ��g�7R��r�a5��K�x�Dz3Vu#&����뭭���`�U���KIو��&�&�`h��/a-�����6��R7q]����u�j 5��>K�nm�,Ϭ���'G/�ٱ�}�t_�y,,`�7�~�{��3!^��ǳ���0�_;q�j���?�ui'��׵����CT��z��r��Y����� ԌOS���aj�Yx��}�R=���}T�����@U�)T��o����M�~O�x�������B�o�p��}�>����.�>���2���h�*�(ɇ��Zp�
M�l�[����Qh?bCߋ_Qo)XT���N��C͟�?/�H��7{�DM��Y��ך��|m�3��&�����;F �6
>)�3P�Y�u�;~3�k�h	)k~J���S�pm~:��3M��&���Z��������w�A�$Bqq�Ǭ�ʤ .�=������gk��=����&����I:��t�ȣ�L�Ø���%��)9�ɿ�^?�����U�6d����DB�8i����)�ϔ��:+`�WY�|U�#/�#P[�k�h�����v�(�Dn8���,ٻ�W�9t��wu���:D4Þ��~Wl*��)��~�~����9f}�� ���v[���AAB&�|A�\Bͤi�c�3"(��������2��u��|J���
aC����&��pL�����	i��������]��R먕X]f/�$�I���o��{cy����[#�$9'�M4�5����hh��$��f,�Ê�e<��ͥy(Y�g�}��n}fV���ď�C�=��[�����"��-}��"��Lz�(F`����_���KҳM����aFw�������?B�odn��b	���zO@�Y&��e�&2��[9�'A�CMd"q��$F�	�����,Nl읩�U����~�8s���f�O�ū6As[�"�{�3�$
h����ե3��A����C� G������5=����k.�;\��u���a;���5�-�^ �0\ø��gU�jFN9%�
)�\�i�u��J^�Kϲe$��&���v`\�5s��j�Ju�_��A�ʵ�v�6E( !�k�\��ݢ�����9ª�q(�1���(��w��+�^t���G�Ep#��E���Z��gY�#����*��ل���.78�HeG�>Sی�\;�<�|�C4���}��z��,�ǣ�����ѹ9a��v66dy����3|�|���:�p��?i�v��D컀�ʿ��}S�[��?K{k�E���1�CтT����T�.BYU�ٜ�b<�>	NZ�Zh��_�h|N�;���3Y�i�LLZ�[��I�]2z��}�� ���xe���Wq\,ؘ�;�~R���f�}�� �46zu�x�d�R!笗f��+r�n$/�I)��6��3Ba����(#A�Q���y`Ck�ջ<��ŶB&��E��� aƔ��tr���uZĄ����
S�X��'v<U�N�jr���^�s�h�����n��H�(���]�rg�_1Hd�����ōe'��<�O�沷d���B�B�O����G�d�g'��CdA#��Dw�/׾��[yL��F���տ���(�S���(��]l���Rm@�k���C ��#�1[����Ò�H=���n*��:�������S��
ј�L*�.�<�x5��>� [�<�����ݍ���M�E��t0V�f%�._%iw�A�:S��g��qs����(����=���HEY>�����J�[���y^4~��������J7�f��Ń����y*
�]b�3c�c�kz5�q�S�	l��K zaD���ا�|�i}^,��x�7���r;�`AHo��DP��E�}���@#����	O0�Ķ�Jif���T�V ��sra�@RgV3�%7jdG���
x6z�t�/�̨��tT�&Gm4�؇����n�R�U��#ZNd������X��ǲ!���U��5Y��o�@Ú0�i8�ӽ�`�׋M9�XF��ql��A�T�hvq��U��Q`q�VClF���evS��N�?���D��ڪ[ʷ4�w?%�&���u������X����h���K��f��0�lI�t_��6��4�&򒌫9�:��IP ���y���p�G�~�@��9�n��(V����R�q�x�� ��P?�_�,��W�(eX��Y�.1=�ޮ �A�L۝�Q��_�����$��1�T�:2���]P��)���/�˃��gVdJ��k�R٢�=R�[������)��jP.��9U��U�} ���۰6����Hq8�ݠv�	[*F�;x�ٱ����r�#�o���[҇ɐ;�����+���0ة��Ż����̉�@�_,��B��Ka�ds�xh��%�1��}�e�y����"5kۅ�ܙ�3;��q)��\��{#A�-]��%��N�2A�*�=���K��Eux�4���u��n�ŭ��H����Mh�>��7�A��46��E��`$/�;�Ɠ�A�Z5�SɎ��t����'�C�y�`�2O�Ϙ��F���` <��u�����G�P7��@�b$�k�UƅҌ�hj��	�t�z����F?���mk%�-���K�ؓ
�P/���V��K�p��Ĉ���/ߩ�+���߃�58�݈y���,�N����S+DKbU�*��f�
�::綤u�&<��6���u_=)ޏ�˜�����ܩ4��$q76@��ÙRR�،��$���yj�E��I�J߫P(���T?�܅\6�����`?���I��7�� ��.G,�2*�g�ЀGߤ?�j��a�٠Οʑ�}[���5�B��!��e���;�{�`)�k?��>�$?��a>�ر�C�Ơ���;Wވ-o�7�
�����+���f����V������Np�f�ͨ�����[�`�yӓ.9nx
�
d��'�g�7�)4$��}("^�����IƔ�q��!�1�b��$�����8�Xq�#�C�Ye��d������Z�Y��SӰ˅�ĝ� 񛻗5H�?l�;8�>�����Q铊����BU Α�FS��X�[_��΅}3�����0���s���f���: �7�k�1�2G��b=_�Z�Dy?6��+�>Qz��B}P.���ґ�U�aĘ��	�X��Eߏ�H84�~���,�����6��w H������d��~����֗�2��zH���Z
�5�K���!��c�Q����0�K�Bi�֙��[)7�Giks�������*��<'.��hS���2�f�}鮿�¬&
��A8y��	v�h/�.�*qZ����Q�+���\D�/D�`C0��-NX�a�9\I�Ͷ��4��}���OK�ѽ+0l��,�'�JyhmP*�q&�=NY��>��&����@K��4Ú<hp��f��\Qf�[���&���XM����ɟ�zu,���Ň�miS�O��hp�E�
��_bRx� �1(�-�nG�m�0"T;�+^� `F�O� 40ɊUXZ��� ��d�M�au}'�Z]�7�em�{���ж�E�E�Kg��\W�eN}:�_�B�&r�w��@oea�٭��֜SSs���G��	5��"�m��U�*����zcQ�6�E�5�E}cGx���L�c��IEjԡ��T���;�i��6���'5�Bvs[�[b����i �
{R9��o+<�\M� m ���'3I2Pi����������n}1��oN���ND�pT_�NN�}-�G/^�ޝQ֎��ل:Û�mʀl���M�%��S"��GtE`�]��S�;���t�l]�����GX�"�����V�L�﹦H�
]
� G���E��2��;���l��*2�?1O���O(\��Ns�+Zv O��'�aA��M�����!ͥ8J��D��.�S��W��Mh�B��)����,�*����+����$��۳֍J�8��ߞӉ�K6#�gX���C�1�D���'���� FOA��'?������g�H��,�%��в�;��ᣀ6(А�qĊ|�y=m��`��R���w�k4�wY.����eqG�|h�S�%$�Gɷ���ʚ��3{���RBn��=�b��@�9;F�+8 ���aKx19�׻rߝ�*=��@`���!��%U���W���]g��D����{�`1`ı�~�-�~,�S��k�=DC]�8u�x�S2�_��T��+�ȹ��u^	�+�I�ܜH"P��� =���J��g�{���#��돬�w�����<9;r����/B�-�!d����=�ፅ�Ye>�X��0�jx��SW�t���x:F��D�1��b#^�{���be�+�9N���&:0�'�\7"�8
��Ȃ8�Hh^ ���%'�op���f��y�
�g3�U2�Xs���hy ��umWGd���ZZX�!^�պ�$�
�X_�7��X��� @B[䖄.8J�'|�4�va�qC���Z��he����xd�=���0���/��8U�(2V.��>D�Z�7��=uY�]u��&e�/�/W(�B;$Z��VCʕd��`}�e�U���[CiL�a��.� �^��o���Khsb�N�H*6ͷjT��' qM,O��]���|�%��9����%d��녹'��e<�`-�Pǭ�l}�t����d��II]+����_�4B��q��"�\I�d��HY\��n�*� ��K��}���r��1	�.��M���9{E���1ƀ�g�&#Eܕ�7��/�����p�|��T�LB.I(���M�oL	���1|r1<tn�ܫi`v$�
�§l���o�$��ү_��,d�+�W�l4��~kHf̢?��>~�3���I7?Ӈ�N����C�$����\���޳�^���Q�e�W�������As\~���Y�\u����n�.4��4�hS��ܐ�x������������_�I$�mU&������Z���&:�!88����}����ڨ�����r�fZ�I�4G�$�M��!��
'��dn#@��L�5j��ױ�J�]��x�б�;��'�$�a�eW���L�(HCG�����8(���h�7��c�_o.�vi����~���u���{gT�2�1�/�j��
�t��-Wl�r�V�\���B����60����E@���ǻ�Z���F�p�yI�TڙIs�W~�x�DX�6�Fĭ2���0��0�F�L50q���'�
�`�4�J�AGv�ju8D���0Jtky^��d3|zs�ڏ�`\p\�<��C�N�df�ȇ� )�@Fg8]�7��zj������[D�x�
8sxS�k�w<f{X�/6�t�h}�<�!�����d,��S�d�Ǩ���e��5l�w���prP����Nu�
�&�H���9ƭs�WGx�4�w����?�;j����XF�w�-�&����g���^����F���*�<��������P�@O�32qjF���IѤz��z�l�)�{%O	E��h��y���|��a^TX<��]������*X�4�L�.���!慙$��~E�] ������\������|����r
CM12��a?���~L0��C�X@䈮�js�ݪ\��(襢�ҖD!��M+�e��R7-U���Uq�l4g�xc��}<a&��"�m9��q?3�eF�/��[�!�h�Y]\56T��S*�]����(x;��{�1��o�T��Mj� �r�A���@G��&,�R&g	%6:�����v�Np����q�� =l:�2C�u�H'0�sF�7�RY���
^��t��u�5�[�1�$��ƞz(�v҃�B��@b�'�9�0� W��;l�A��A�}&Q�����O�9tv#%ב�@ٿ�S�C{#=V,v�}䓾Sx;�2y�ܸf���VC��B���ʰ��!��N��_�|}\o�����P�;�D���a�"%�wv��˕���<A[�{%�}��.�`�m;Kn��rf����^�D����E��)��>��Q��M�Ur��C��",T������+��"��l�����R	�5�S�(�QO}섢Q�Q���Zݳnc(�q�X��<P�r49&���N�*�E<���	AO�UtO�c�]��j~UcY��A� y�Y(��E����)��W
d�iN=�y9���ʰ�5���CZN�w}��E}��(�+v�f�J���f��H�\��$ޖ  �}����`ٌ(�a�E�%@;��O���#_ޮ����cɴ���\�`���g�l�h�Z'K���U5���8�0��f���G綪�vR���RL�ߴz��`h����������}����~��3Υ��i��9Tu���h���jq)����Q4ᗥ�T�OM*ٴo���<���yf��9eU�����ũv�7����QQ�%�b���SQV����p5�ps�f�N	��cL�7���`f��!�r�KCe%M���=A�(��,N�ZO���R����귛S5�?�ԧ̄�P��J� �*�]^1��"����؟Z��@�&K��}�Ɵ����i�F��B��#�ehE�l:����βgX���?:'_�N�ڒz��'h�l����;��Z�۷�ߥ��������I�X��a�Z��\���DK�Q��/45���rD�Q���&���NAڌ��0�fBI�m0j��ov��$�C$mR+BM��&XW�RP�e8�9��/��ҳ������3Q��p�˽~�b�<�rU�ɮq������\<Έ|t7��&��`SN/Xr�Ƚ�V��ݳmfagd[}���%�� ��k�ҏ��G�iE�Tg�4ܵ�b���Fד=#Y���'���=<Jm}���Fr=[7P��I*���^�#���>@K9^�u��
W� w��*w[�2�^�2����w�/�����х�A�޺eK��>%)�X��o$b/-ZE������|=��e֦�Q|�E��&�R:�Y1&�o��MD�}/o(�@�T��C'�L�0So�Lq����Nr��F\�J;�zzyd��x���ai9!f^���{���h{�:�+x������8�4����勌ix{`	�)ca�Ɇ5�����!�������������+��AE��[I��PlA��R��-���F=�,�ϗ�t���/�U1���_�w�
�����Q�����M�}c��R�������M�J�s�����'�HL܌�����?X�20a)�/%|���h�7"^T�Z,�x_�xz�3���i8S'sK��G�鲛?`_6�JZ-*�c�I�`����Y�	��ҳ�Z
�'!4SH2���:��JY�`�O����}~�H� )��tw�ͅف��oa�RŖh-ǀ��]�t��4��2ԫg�c�).�N`��~%�A�oO����$lx>��1=E�����t�����S�AG�`�9����?�L�Ӕ�ΪȁU�X�>��8CQ5t�Z�;����#?I����@�\���6��p�e�ڍ��P ���H@	S޴Q�D��Ҏ��j���X{8�Fs�S���FVg��ބ�7����g�'?�]BD(~kvj�
`�z��#Q�¢~m,1��]D�=����lu�������r@��s}*	;�⦅�K�)c�l��>>��oa��X����ܓ��Z�SD�7w{U�2�ܑ(T<������
x!�H �L�f�ʋ�Tv�Xh%�f���k,I3	��'���@�u��$�[�Z߾��酕���#e�p{�V�l@m�g�ƕ���,��^@����E�����/Ϟ���5{h��c$3�\,�6�lL>`e�s�6/O)� ��J;��1�`n�#h~X��j�l.x�
y� ��C�#�m�H�a�%;J��v���$��т_���{i�<������̋Ŕ����@1�<T5��e�T�ȑ7����OZԙ���J#XE�YM	!GX��niq�eY{���z�'��~�?z�`�'�іI�$_�w��+[pW���������D	~��H��-8D����$|x!>m��j��=j�m�k���k[�Ѽ�e�?%V[Y_ٮ���5P���$�"f%�q�M;������
wԿ�h����#��n5���<�hq��'�lM��֥���=��{ ��X��&;�	<QQ������$ә�2�tg�8�K�l�J��n ��U�>�ҡ�vN[�(�M�����y S2���^�8��?��Tc<&�7joͦ��H����9&n�k���c�e�ZL�,X}�%�	X����S*�FuM��6_�]��8��8����凛�}G���<@x���A�:Vz��Cg�z���1�Z�2�!�H:���Z�^N�Fj_�Nc��¥��d��e R�sn��8O��Cg���$�So��<���|����"h�S�
��S�V���ƻ���� �`6;a=z	R�жp�#����E���G�EI���xԡ&���=1�{��h��Eۄ!�*	�G/,u3fO����ݢ�BNC�4�2��3+TJ{����&(vu�6���z&��_��G��S������FN*�ؽ�R�A��A1�`i����̜�o��V�sOx����J��(���ܫ,��s��O�d0d��9/��� ���P�5����-曲o���ʂ`P���1�|H8	<m��t��O/ed����f����i�������b�<��H��c|=^��߀[,���`��°�+�{��-d�8�����ܝ�0s�z������3&|
�ͷ�HG9O�;g��n������ŷ�̜v���j�����C��f-wS�C��h�K[�P�Y|;�t�����KSN[�� E77Bp?41pp�>���-����Иx��ڦqx�o�
2� �A�@�!C����6��G�u\sH�$��簅��'�A؟.4�I��8��!o3��Ŧ����b�g.�!��	� ����|vC�^b��)#*)䣧l-BA_M������E��Lg��@�C�ʌ)K$0>�a��xM���>|�`��/�s��Z��k@	�Sct������>�4���/L�E�s�:�N)'���=g�@��<$õTK���� �'����i�Y	5�L��@(sm�E�������qZ�U�/k�[�D�Y˧�G�ʷ�y?J����DH�=j�]����@7D�J´h��0�}��n�M#.�q��2=��|�J"8A�������<�Z$��g�|�!Z�anM ������y�gǮY«g_��4�sN���[�0�� t�sDi`�����8�E��-*Fyd�� $�;֏��)ޛ���G��]�5j��h7�(�*O�������X@!�;�fS?4�Ѹ��Ȩ1�}���kU��C�g�yZ�����(Hf0�a��n��2����ap���� +:u�-�����R/fa~*����3l8\���no�3�R�GU��	��5�i
�!�-N��$�T��M�_o��|�G�m�c'�}�4fc�;�]����&a�O�v3��>��Zgգ���֒�aL1��͋	 u9��1��ݛ�b��.�҈$9�8�����0*�QU?��K@��˳GVV?���Wi)F�c�;I&X�&N%{�}k��O6��R 2�ԢR�/����o\��\���\C�q�M�ݫ��Tԫ�U��(�&<j�)D�(�TCG	���VȚ���%b�x�K�F�`fQ����4���������ve_
�͡,ö��%?æ:k��u���-�S8H$�����b'Z��g�<mGRkP�MP6ơ��;Ia��������
|,
�K��E�'~2���7��,P�����:�=����`2)��k���%�f���.�l��/�vo��҉���t	�)���A�Uh��X�N��PLV^S��n���V�i���dx��/�4`�μ�D~�d�� 3s,��p�H�q�ҭ(�����ht��5��
�d�_�v5E���5���C�tK���)^���Z&��ï*ZVK�gϩ� ��ꯔ)�F�q](�����v����;���b��w$�,����=�xfF3(�AE0y�L5/�i"�)������ݩaQc 
uC�R!�_~|���
R��vX�e�T �~��[�,;��Ht4�q�ܹК�,o�I��V��l˲ߚT!���Q@����.ء�t�%� ޶��*x�Oz:k�!5�A��cf�/|���~5�C{�]#aZ|:(�5��|��[���Y.h%��0��{�@�]����W��V�`y��pH�� �|'�G�rD�frǮ��b�i&�I������0|k��=�e{��dEI�I�!�c�h���l�7����-�������4'�v�a�|,:�YY���ٷ:�}FT(X��1����&e8f~d�R���c�?)~����XS�f�)0��ߕ�ݡY!BS��3ϔ��$q��û祼��Snd���U4�?y�]L!�P~��mY3d����SE�`�,��#��,�����GG�c���/��v��FN��5V�u��@���vW�;\�8�9�����}R_�e	e#%�Ǭ�+���w��m������d�ݧfS_��j�[���A�ˎ��z�E�a�F��a'b�:'�OɎ���1�3De4��|�+��V�5��N��Pjf$'KEC����s���nvp-Y������3,���Ɇ�.�4Z���P��v�E�m�_�s��z�"�ۂ�Y ��.�Ql�ov�����qtf���S���M��U�n��'v�yZ�i��-@%�&�&�0�־�⩏i�R��OnD����`�ii$ډ���*@���c���X�G�.yk:[=�>.��ޖ��aG�tD����6 �\�?��6�P ���W�Ma���#�7��o7��[!Ib���̒�7�,{a�\H�����*�=!x`y���@y�_���*���n��&��]�aND�F`�������<q>�g�-^��-�/�l��ș�ޞ)8< ��7�B��qs�XEm)�b# SDe������U�l�'>0�@-#� �͢�}ڊk�H)	�}�O[�ʱA-u��]Ҵ�~�b��_�,gڼPI�E��i��┣x�T�I:X���2y��Cp�ET�B�f���3'�R����+��~S��2�����'�5�*�Z'+_�5��(o�h{8]K5,��PuII�je��-o��iK���8�z��"�]�����5��UZa��!��=�
ˊ��y~KttboI�p|���>S��K]u��d�>9��=���)E�W���[ܾ�Om������9�(N������i{����#y�ɗT�V���x7����?���2�(d8�W�=]@r	�Q ςl��2<��XxKu�ݙ�v�5�.�1���2�]	t��
3{5|_�m}����p�a�c� �<���YBN��P���o�!P������S%���s�L_l �p2 rɘ�	�V#�`	�����H�����\- b���"��e���#�X;Ɇ���M��*kj}k�B�PxX
U,����"��_Q��	��p=�T��x��$k���䭦qh�BPP��P0�/��w�D���"�{��� �5�M�b��H��R�C`��
�A�C��r�[����Ç�	'z�2EǤ��s�z)���7��$1��`���T<�^o}���.��v�1��"WwY6m��"���ͮX����P��a��R�v{|t��!M/���F�8�&��a��������K������C��+���M#O��& �3���g�30L�-$�������=~�E"����	5t ��7�[n��Oy�	ciNaS���@|���'EC�D�G1װy̤��0Bs����ԍ�q|�5�r���m¹�gB�@�z��^����j8�4�T;�lp������&��$�/�u��/@P����>��Щ������0�&�N�ՉX���k�H��x�iYE���*�@e�f���(b%,U�v���NCR�dd�#���khx�z֓^�hJ�ퟪ�GK�"�Oq�}^ȉM��\�dJ�X��������;�
c����-e �'��1/!=�?[3C��U��w�:t�2,	y�MQ�?���j����®7i�O�Z�^+U�/_���t7}���ŕһS��#q�)�����	5�(D/�x�����(�DϾ�"j�&����,�&��ah���0e󚭤��=���V��C�2�#17ޫ�M��f�4˶	���!��;}��\�*�opI\�HП�O��JrN>���/�B��
���)\�v,��V��Kz�(���04����¶�f�o�U����y� dؾ��q s翗l���Y�rZI�!|Rϰ����bl����eyE쎑�_�+�����%�٨ا7G�Y�R�r��D���;-�}��߽��'1��x���
7� �2.���t#pf�WU�s���Һg��X$qcDg�&^�2��tc�^˗D�K�uH�O�l� PQ����>Ϝ���"?e�ī�L������ՙ������JRcZ�d:�Im�Չ��n˼��P�����r4���)��6���h�ZNy�ls\�|��� �ǩ��	G�jU�&\�j��k�����ʠud�$S-6��ݳPK�ը�SF�D)��Q�e�R��s�8�h,��n��������~����z j&�����B���W����L,��ফ��E�Qu��ι5u�,f�o���a�ʩ���|�y�����@��c�tG�P8�$Rc�t!I>�z����\s:����:ob&�`i9�im���u�c���fN#�1���X�UIS@K�u"w]J�b���DeΚxI{@U`0��\�å��_�b���E�Nv.��F���-�=�ː�j������z���VgƆ�h9�w�!�����u��$WIq5q��n�/���K7j���dq׏<���N_6ɼ��*�A��u�Iȶ�<�D������}�@3a�b�B���#z��3^��� �{���O_�5��X�+~	�eA*ť���P����
z��zK_��R�&��@�k�����|=o�����>Ei��Z�[?V&i�ݍx�<��g���"DD�*W���(9�@������H��p��qz�u�]K�6�z��	��,�y�}k"�紬����o:��M��)���5��'���L�O3^3Wq-����,�8>/��ka�&���<3��N�L�M�&�4/��f�&�d��1r��13_%@8�oOpr�Y���Q�(�D�Z��*9�(p�jTRձ����`�.;�{�_�?�Q��|=|��ݠj�Y.}�+RJ����GX��_52�4B/l��raR��c��U��	#�:N�Iy:7#�D#]��Eg��wɰ\�Y��[�6!e��Dn�����Lj�$��*}�)	�S������=W�	�m�B�[�zAp7�|u�-�ݝ�i4��><[`���[���97�Ƅ�G+&�������%��-}�[{�A㜄��؟�{�$��8OKH��'�ΠB�����nU���mXNyk����Il�P�$�i?>|3^e<�[ ��;s��lrL'L�����m�
'a�#����!B��
�p�����=I7�>n�S0}���>�p��(��|����\���9�5�#f����`�x�?|L��������xw��W��HEJ��������=��d���$�C� �l�I�іϕ=�:��ڃ��B	S��ux��4��]8|?���w��*����S�~��4H"`�dǇ�{���ϙո�c�O$(�f.�^�<a�+q��ȳm.h���]DK�ؚ�i��C�BϪYː֚�Y`M���Z<#�,p�eu2��W�����t�a{/����[.�M!B��M�5?4ض��] o[-�S���19� ��GWo��@�2E�n�D�0:�!&0CO�7�����iñȵ��F��W�:1t��6N���^�QD��o�Ɣ��Jj��fg��n���! �"D�7� i�ڵU����,��*OV�$<� �u���ׇ�P�Z_���R|�_�'i ��e��-�c"̏H�r?�|6�95TD��J`�0��̮m�w�lf�����u�^� �,��x����%�!#F���� ��:m��X'�]1�k�֎4���V,�zH�%e1\M��J����Q�'����l��扴�a~g^�jL��^�?�_�Ș-	���Д��?K�.r��M}v2�Ӊ� D'�2�t�o`��9{ٌ:^}'%'%���J��
VA�Hg�ƿMr�I�*�K���+�{��ȉ4ɏ�;�P���Y̜s�'{�	��ِ�ԝ�̤i!�}���tѽ\{ބ6��5T(l�e]b�\!�4Ǣ������-IV5��)_���}�ߏli�Ŧ�M�d>D�G��l���R��6�z�<��D�Ų+4�
��>��f�C'����o��>�"X,��/�|�ը���d�W�.#<�E�d�����q��^��N9��@t��cr������2�u�h����?�8��fg�8/,ч�����zT�KE��Y*Ee�`��#��~��k��)�����<��[�m�Q��_�u��0oI�!�MɸZ�Ӱ&��#���"OP�Y���C*�J���N��c����4Ǥ	־�A#*�"��L+���nZ�Lz��N4�l;��|�R�@�=�4�
���`�\�e��� T[�7%9��2���p�\��J��k�hSC��b���g�
[i���.!6 ��]�i�5��a�	�I�o�%9���g�CW�0�Wz��W����*^�"��W����gs����}\IMA%��J��[!�1H/$�����}^��lB*�>�Vq�bcA��b[un�d0�_4h�j���}���7����D][ջ���,u��t�����bΏ�ЂU�D���������w���5-����А��]��{�5�5K�+'��5�����"T�x�j�Ym�ڦ�q��v$�4�����k|x=�hrZ�/ K���?��M;�՝�%��2�W]�9t>�����k{p�Aq���z:N�\�"�"zM`�����;j�^Q�f~/ z��� �S�ў^b�7�@�c��
n����1��'g����u�G\_���W�����wL�d������hϒ�6 �������~%��g�f@���=?2nY|q���#�JU�Lc%c l�/��r'SN9�b{�y�?�
B��[�\�!=1:A�G�Z|�z��^��x�q�S������ϡ��L^r��fB�
��j���ɛOB��+�/�1�J@��K�G�`��
S#dك���m�tsݹ���!��g ��7�x�!�ۿ6��\��Cl�����<MhO���xZe�u-�S��uU�9T�耑�cPRa���ǭmA���z������ƣN��%%��fX�5�K'�TO� iw�BC�ȿn-� R�AZ
�:�������������ho��E#Q�ž���F����@w�Cl$\� �;CY�V�[~�o2���C�Y+�^��GV.���T�<i�T:��ҥ�������Lm�&�%~gC������n�a���i6M����"�?-os����iR����3�
������tPf��Z�N�-��S��s�O���L~+iX�r�80����!Pr�a�V�-#�2	uj��`�(��A0���*���#穰�붆t�_v�Zv��3X�6;|����K<M)����O�K�Dţ�Z'Jf��U3��9��(����l�2�vXH���s��}ߏdo8n`V��mk2V/d�A�������.8�x�l?A�O%oJ�"��8��}��Z�97Z
�7Sd9;�٬���d��35��B�u��D�	�6�T��?g.��sM������j�A�!U�F���a\� VH���0�A㰺ݥ��nW���~s�.��JY��#����2Bq��w9S�g�!f�$℁_�������Ԥ9hW��#�Y��/@�8m��ϖ�U_�|X���@�<�ؖDRl$A?*�~Ƅ�ҋ���{^�n 
j߃=%Ŭ̆�fg��C ��UI����;�V�x
�ŝ�;F�R�-�M�!�u3���6&�f�ȕG��	c�O���2"�Q-���>A��������*z��c
�'|,�x�$�n(���jx�δ�bCgܗ��"�z��-|S�5-���i������Ll���Ub�NsC	�>�A�[۩b�S$q�l-��E}/mgQ\�l�����	��D�P�S� �~�FRUu2�ṀP��gI� zA��+'�8rt�4e�կ�@��дI����rռ�痖�j�U���n`�=��_��̇��q���E)� ^J�86>@��g�t7�9 �cxòb��m���r?���n�J�K��C	\[ז%̕�N�����A!�o��u���}���_Tқ]�2/�SU�5E�x_(�)z>�O��oQ�\Hּ�]����Vu3��lAጫ�[�.$\�)��T�4-0��g�������-`}a|����Ǟ�{��iT0*G�l� ʬ�i�q	����~?��-D��q/��M��}
������Hϻ%�[�-M�!�i'��c��.�����.w��,���ˬ�����t�<�[��@����G�]R�6��ٓ!�s��$�w��՚+�w9��)�{�)��rUZ������)�}�Ѥ<�� {u���@�|�^�{S5mSH��~�����������&��P���D��Q���R�����f��T�3�l�q�j���Ggg<is��u+ܩB������shsD�O���� ٔ�� �Dmk�<���:^u�[�hI'��r�͍YX�8��{�L�{��n׫��bH�2�Y1ꔣ���)f����9����Z��Du���2k^N���$
�,\���UO��x8�?5�ߵs��yRi�c��p?b���uU��q��h��y��,�%?�jZ�6��=?MB�`���������t���_���@D x��[��Z�m'5�w�����`*����T�6���sa�g(��a�/pR��T9�u������X�?XGG�H��)�����Ò���q���NdIc�[�֢6���Ұ&k&�l!�o�VlHϥ����1�~�ˉ�8O��F����Eg���`��>���ؤܿ�iS�
������U�8ʎ�[��}�m����́\V��z��돮���}1�� ���5 ��
��9~��l_�L���z���mZG��l�lʆ��"� Q�_-@}�+�L� QY.�"*%�M�4+����̬���.����~8��d�q��\��n��Uv�IARQ�#�
� \J��y���J�3P�E&�',���"xxA7/�O�;�7�ם���*<3���ս�,x��ٲ�T�Կ�5�R����dkx��z)QF��,�K��	i=�Ц����_������e�Z�`_��@�;�#y���:�D�0Wd]�IEƜ�4�H��ȾTėT�b߭��(��z��^��g7�dg���}]0��}���`�����5Oh6Me<�x������c=�7�""�݀��|��݃�4���/��c�!â�K#\�.詇���`v�R�y((T0�-e�Z�b� ���<f���c�;��E�&b�R:}ZD&yC��x���9��?�Az[��F��}���2LpFz��r� 97�ǘ�AE���W�nF�
]�}�c��u��=�9e!���?G���ŋ��A�9ٺ�t�o��%�O��{�^��ƢЖ�f�fenN
�i鍡�T���rl�0�
i�M�"�����hK��H�	����B&z��J4gR2�ceF7�=�z�_%� ��=!�g��p-V�&����=��w7cd�HyN4>L������v`��.���r[_��=��T��dK�n��ܝ4j vI�`�ܷQиF���L綛8{�c�Ѯ1�]8���M���:���D���dT��Z������8�Z&�-�P�+\~�SW�j��T�-��'�	��8��^��y�Ӝ7\_��3JؙA1ps9�����4U�_��b��W|��v����~R�2��^
[6��j,�/A���~e�j�C��2�QT�h���	���T�ܷ@K�����"������L�g	�5������#4�>3D�g,o{��xER�nz}�e$4y�r�S�t�5����c��A]������#'8KU�0�:�q��jj&s�Ԛ^����:�Qc_w4�G��2"�߿�
�)F��q�Fk,1i�=��?�����=c�Z��-GN��=nof �~�o���ʄr
I���{����ԕ>��|1����ky���@9!5 q���`�~!�{�x�����o���mF6��γ�|F%�ۜ5w_��n����Ub��_�B���m����~�'�̤i��5���b�t��e�,ԠiB�YXZ������`~�G��Z�s�j�cN��AM��	���8�AA	I?�JC�v!���{�a@?\�pK��:��;8�y�
�a��Ǡ�tCՒ�� ��B���U所`$}jE,Ǒ��R�!�2������V�>[I�;�T�'E1+|��\H��ΰ��Ŝ��+����S2�p�k���/<�R�)H�Y��qNW[PHI��(��5��ߞ�A���������/vޒ���'�v�?E�L��?X����Dkp����t^�W>G��r��g���L���  e�/�V�d��6��r��Ppq�F�4�|�>W��3�c�]�Y���q�D�y�ǦK�¤4(���o�&-h��J�����h�h���3~��Bᒚ� �0|�����>�C얤�X��XL�6�S��9������j^tu�M�a���
���EBܻ�����%����R�1Z���"?�&���T��iE��\
[+�=���p�p�O�;�Βk�3�^Ye0�h�#)M���m+>��c��2 ��M��F�c��'f�������tܾm;9	���N5�4��p$�25�2�t��8����t�]��@��g�[wf����NC���ԀǙ	Gl=�:M9�R�,%y�2eZ�����<ҙ��M e9b����#���Vu:I�`M��a��K56��R!ˁN�"�%�C�Cڰp��5P^��&2?�Mu���/�m���S+S� a��H$f�_d��l�C*�NܳWc�
__E�����Tͺ�ƀ��`���q�?�"[���t&��Vs3�̠���$�͢kIX_�4��L}v�]������-@"��P
�(͜l1G����a7����j�&륍�|����Y��;�����ܺ$/k/ �8�fq0��OW�6��!��"�kh�<vC޳����@���s��y[9���ۭ�.>C���?ҍ3��L��E��K�_�����-�S��߈�J�s��V�'���٭�g�]�$�(�H+��B����^��z��HLX��
��h����U"d�;>�~�p^P
plk�ϟۢ�x�M2��#�[� d�k�j&F��6Zm�V����h�_U]��_������m.����ܴs&�����c(epP�����[�P�(HK����s\���;��	]����2l����̲`/�6:IA��~D\���pk���=�Eh&s5� ǈOq�����n���4~9U3�9��(�1�f0�E��,C��Vuvx-����Nw!r��|��-�?��W�J6�+y��?��ΐ+�;Y�M����� m�yJ�iq6�+_�n��F�-�>1��̞sK��[/�	};e���cc�-���)���1\����tg��\>K�����rm/��{%3�͞�������#�������}
J�� Œ�X���M�5B�t�ϭ��ƟkV)(��F)��X��Y �_\{i�p�Qܰ��?F4�fE�Ymv`�>�s�!���4��H�,bv{广�D�Y����h��3�B��;L�[�oq�.>�X| �����/�(������hHbq�[b? .:��SQ؁]JF�e�a��펯�O�#�����<y=A�E�x��|��@�4���E��=���1������Q�t�/�?��Z0s7]?�Ќ��%�U�1��M�zQ��(DgPnbX��w�)�z�X�7my1�
Y�!1߱K�PnW&�@&�����t��1����O�]h2���%ʆ�.��ǰ\�XM�˹qm��UXt ��`�/���:+J�aT�|P��3xM�#�M��m�M�滙m�W��t�xc��Up��p4��qx�� cy�?zvp�I�]���UXt#$�iR#OB�����9x.�Ľ�@ x�H3^�%��}�ʍv$���]����X���&=u?��_����Ƃ���Zԙ1ϯQ5K,���F�,�&�?EF��ˏ6À�V!r�t|f����v|J�uSU)FR����C��D䡡Me��}#6)��n��@��z�?�4J��V�\/��a/�ԥ��oJ�?���͇U�����Z��e��=$C�~�.:c�E|t�o�>J!C�1K��(�&#�F�0P<eI�f��fXV��7>�^?��7n�|����C+(xrO���DY�5j�<@ i8����8��[�q��I���������ɛ�_���&G���H�q����A蹬))�����~�	�;W��P�B�����>k�3zt1��B��8T��i�9�bڅ�ޔH	�;�I�Q��d`8/����r��w�"�'�#0��%��/iC�^(���}H�f�>o��-|��Rk#ѡ$��=;�:I�Ӻ�edQ���t��3mi��H_e֙�STb(��-gI�
`�����4%��,�)b��#N�}���i�R�j��v��XVb�`jYFŲNt=nE�+�%BLs��lN U%����]ZEHҭ^Y�h�����ʸ�Vp~BW4��qr�����ĩ1ym�i��^t&O\�n����&���^��U�>a���V�q)����ν2'6�r���ؘP�zO�;SnCi����M/U��]�O��08�趎�=��8��cf_q�����|�d[�pDf ��%�ԃ����3n��{I���w�r�	TU�b�y��`-F�Q��E_T�,�%����)�
Zc�.��0�����P�yX2J��Z�-z��d�� �\�u�Y(i��,��Դ�?Y�2G�GG]QQT�6�`�w�1?���6{�	Ya���+W�R�hd��Y�mN���T �j���KQ_��-U��^r7� !P,�@e����ne����>k���㺸�e��� f�u{�ӳtmW�@ǕdM��F2͢����~^�8~��@`�gso��N ��"�n^)���P�`�o�FePa#��)�$�V%l)���*��;�@�R<΋��`���h�f�"��j���j�Т���lQ�د��:�^�"5��\�dw6K����j!(d���a�K�&���l���5~4���n�hD����[�@��k1|����8z�s�#�]�*T}
� ��������qY*�O�R��C>P�-Ac��bf��,Q�_��(��	�u"��nAt�&�/�;�����є~w+A7�E�[6���$�����2�'J�N��`hX8��u@�uUǧ�������4�����^�8��`�K�wH �z�Խ�S�F�u�{lx�]=8�X�BS aFuUy�ü$��qG�(!�$��@��;@ZHƏ�$�,SgL��תKq���\B�N���/ћ�N�j9(t7�b
������S�;��J�hkN��3�B(-�AȈa4��L�$��<��K	 /z�tN�v��GV:��p��>��y�[��L�K��P�y	�x,e�W��U���%e�/(�"_T��4hg����eb{���?�0	������&�Z��S���`s��5Y/��'��M�~��3��.c�/�����b�&  ����nb=<�y�S�+`�t%�ATG��}���^��
�����ʣ;og��A$��6��hj�(1\9�f������������^���Y5gYG5Ӽ��2�b2Q%ބ��aCvr�k�*9Qd�s� �] L�^��X|�z{�z�`��!���9���|@=��Tuc�_@�ы:d�|t����"fB���Xo���s�=p]�s�F�x�n���f���͝7(�_�!��L%OV�%8N5}�֦��7��4�B���Y1�f�����O�q�9�|$��k|��@���p�j�K�g��b�H�2��ҹ9��-�L��	��5��])�������δ��$: �`�7OMЂu�O�����1x��tݨ�����H��{�V�r�#�6�	��?Ӳ����Z��W�m�3���M싨�ѱ���jǄ2)D�dt��wQ�?��rG4�hf����A���~�6_�'N���U��l�v8ͬ����M�
�n�UN�@�����M����rI-�#%b�IV�����>�os	��"	4D�x��c������o/��}zb.��q��Kۀ�l
��"Z;(Cc���e8*/O��$�v��x��a�+ܫ�����@0�M)�6;[e ���cc"���5lu��l�����H��:�9��@k�jׅ�X�/���@�3W�(��i�APǑ���ҪF��Y���v4b�Ix�H~�����{	��d�M��^�Д�ط�ea�L�ʙ��۞���ϪL����}O+M�`³���l/XYl�p�o��b1LN��Bn偅m
4���0�N�Pv�h8Ie�B-��%M)�n4��0lV��f�����E`�j��l���6���ԗ��Wg�	�I��49��WR�moD�g�@�;a��C�}��0�t�^
.�l��n������r/��ح��^���;��?�b
��o߃K$��4&�E�7�L��[?�cJM�٥��
���w���^��<�i|P��;���u�$PM�	+g�c�A���&�
�uy0���u��^��ʻ���^���	�#{ϳ���	l�oS)�"����gR^��g�9�����H1��t#~Eq�\%�!�\
h�#�d����!��|��+��qŃ��:$C`,�*���SRD�X���&���& ����p�.���Z��ܱ�8p���=�F}D'רа(rD��Jˤ�Pݥ��"���D"� �ɭ�o0 �w���.��'�C�e��Z;rfHU��l���g�ع�!?�_�!��ɢ������]3X�e>��+��
]�:��D���)9�bxD�����R]���O G8���&�_'�-�T_��J����Q�g�Nb�Pm�������}�)hbw�8,��@�Jg�eb�	�ILbP�Z넝0֜y�J�'��<Z�z��E�qk���yir���5i�œ��r��bϯk�����N0Ã����tX����S+P��s�$"��{`*�ϞI���`7>a+쓌8�g�����d:X���WE���t�]�r��/�zfߩv0��+Uy-��2�e����a�57	�w�5���G�u����DS|^���T�=��M�n�e@u�5��.�-%`/C��r�{��K���p?��O�F,d��0#���kP���I�zV�-�Z3���م)�������}�	�Zθ��5�}���M�V����^��"���U6�Zw����^=D��BA��FV��U��7�ϭ�F�b�o��/�s�qh��2!��!�?u�.���Ƴk�H����ߣ^�4\KN|�����'�C��2?'�h�����ͫ�{{��L,MXgNt�Z3�!d�x�V��V;�h`�fd��kk^��������cI���po��;9��/,�l���!Ы�s��.f�+M�Se�ߖҫ�!#Q�����y�������N?l-?�țgH�_���JUd�;�X�sE�L�bXwoϴ�+ "�]��/3�˗�Ύ��ơ��ޝ�eX7��i��.���&z��.Wҏ��|���rጔ���%~)j<ERX��~�-�I�1����8��2O�x \�u��9)��2�������{���i���]���ea��Zd���i:P�'5��!����Ǻ�1s��]�3�}�p5�s�YX�&�6S���D���m,�`E��u��t�yC��L�򐅍'9Β�4f��Lq=�*���,��&�x4&Ԋ���YN���[W�G�G��c�P?��Kk
飭�@'xu�z�
8[�n$�_a�̩�E��$k��z;�h�ӷ�(7l�U��A%6�_��������G�!�[;����n$��t���c,��T{��@����'|�8���*�	��%�xZ������L𛰻=�t?��]�B`���>�(o�0���΂'L.n�M�(~�!)��P���x䴡K�}U����2� �H��ı���V��>htRڬ�&h;r	�X���K��o�^�o�غ�3r���vQX�$���u� g����|��,�}`ě
)���epvs��x��txG�J�>�#n���2��]���;5��g�+}�.f� ��:�k~�ɇ/NY�JA'1M��8�M�X3C� }u�c��?<FV�%t�fG�M��$�~� �8������\������/������[kӨ"?�tW���a���jX#%�	���3�|$yݚ�������%�H�5�r�O��33sT�k ���ڂD�Y�ܜG�FF���h�n@V���W�˾�t�}�Z�RT��s�?�K��G���hk� .r�x��2^\�T������ˡ�B蠬[M��G:DBv�
��Ą��kj� �.����6c#�U�������g��_I���/,݊���FW�EڔG���̌��ǂ����"��f��#���"��_(���C�C�+g��% x�L��tE�4*��Q�Ϙʏv��p'dox]/V;ed�+���z�}G"�s��Vvh��G���cm��郋��_��:�pv�v/��_�h��H?�������L���F"ԟ���2c-x�;�9�2���m>��Ɵϼ�g��H��gË+3~��4_{J�D)�m"E���uF���,G�$�c����
[ZB��ݚ�-"�g�zp���e����#�3|��_
��I�Xg�x�9 7�i�HjꭚM���z{�(��ؤ��Rc�_��yFw����$�E	�_�$B�˚��imt��Mn�}ޕt�F����&+<t���G����W	�&���h|���=;�OsD�D�^l�QAl��k�r�x/0��v-˚��� ����gp�%P�5s�i�zK��������[s�Ew�d�AL��A@��I��{�^�[^o�r7X���0�ܷ�7?��_�[������L3�t�J�b���BRFH@�(�]�g[�B�5��~���f�1��~��E7��jJ�}� }[�آ=���>�쾧0�(j�Ar�D�v���\w��&ұ���5���(?��qAi����.C+�fIQ�<���W��='{S�:o�(:&�=��d�w��M�WX��mN��^W�"�B�Q_��H���HN�U�ue?o��%~u�֏�8�fy]�~���g9��o��-�6SF5�����Đg�eJ���7�
!�N���u�[��`������2k�ri�ˌU����i��(��{��>\XP�=Q�Qd����u�\��(7�-�V��.۰�TdQ��4o���Q��2���C��"�Q��VX�L�W�vK���r����φ�@��++`s��Fn� ��K_RN)�5�O�C��̣��[�>e�&��36]�n_��e�p[��=�s�5���y��h��llp�z���W��gLm�8<K,�)P�0,��@��q�� g��U*9N���	�3�彘�qk�L�Fw��1dtO��齨��.��?�π8S=�������<��@(���Gcr�C��'FD�T-��7�3�
I��=�B�����0z\�8Yi�V�/4��)�E��{Q�[3��F�rZ�����.�(�$������i�2re���ga�`���#%�0��c�-���w3:�XFIb4����M�f�/���Y�4bi���*ES}5�05k���y��KEU��V�u���h�y��o�G{Ff��T�`
� *��m�{��C�Ա:��%��x�}N�#F�B�$J�i2p�_����HUJk`u>�kst�T�H�q�E�N���DPhn!v���%�5�͏F��Q�� ��ݝ�s
z[\����/��om9QŊ�z7�zWC~j��y�cI���ȵ��P�W$�g�"���p=�A����J-a�>�3��%��!�3�h=3�s�>i�$m����K|�S�BS_ii��`-�����B���OH;������4ʊ��f�����s���~�=ЩNP��[��.̑kk �J�ѯ�FeJ�)�}�=ڐ��g�����u��������(��2�94n�pQ�����y�{�yE�;�%=��P3�WBdڳd�#�@7�V��Z�
\��̘���xT_-�ы#{�����jjs�?��c���da%`��=���ʥM��w�ӬĖ�\��#����z�GrLk�^"�s��W~�C����Ur$���ؓ�x=�C��K�榸�W����b�Ic)N�Lt�yҺ���R,��"��G�9/�ą�Na�.ƻ�]��+��~����aT_�Y���̊ׯ��OZ:�����}N�֔�Qݲ�5�Z!j(`�Ze�����1l�~��`�[;慛���L��N0�i��9zՖe^ҡ&�G�W�}�S��dҡ���F�'a9Θ�6� 1vA�U��rf[��{YHB���+ W;7�L
��z��ב���9q¿�aj��ͺrؒ����� �c���!`vq4-e�#�b�mxZ�� 6�5 ,�ə4J�����[�b�Qo�@x����Tƪ����o�q��%Ⳓi��x�t����Y�LT�ݵ�^��k�Yw��p�{3�}s �z��O{d��;�@	�{�}U�5���j䙟��Nh?0�%`f�E�B�O:lʭfq�}��F�ne��-�">�@3����H�E�L�aχ~����Y'���eV�e._�b�.ibV����$ԍ�A��ɀ���#&�ɒ*�=�5���K�3[�{k����(�����a�vya�a��Y��a����b�G�v���$:��խ��)��M�q�1/��%�o�~�N��jP�q�pG�8���(��-=|L��5�T��<��\�R2�����yLf�r��}�1�]�Њ�)I���,��R�N1`�@���
��A���Gn�k��_8�N~tT5p����a��dFn��W=ٸ�}M��� 7��eP��Is)c�`(-@��AtSG���_±��"g�2j��ȣ���w�5`�Y-O;[����T�/��%���L�B�DX��T�����I��:����;�'�jF�ߝ�u��W�S��C�zշ������<g�e�K@]/ˉ)��{�b�Y��]`b�!��$�\�GS��p�e��-��Cc�*�jn8�D�]��c�Of��C�[/���4?�J�אIқ��&��؅<�3]Y�y�������l%��	$�p���������UNL߼���X�%������Y���S�!�J|�]����Y���14@�I��d_���#m�R<���{��0���qW�WxP]z�p�t�/��߹��rC���/4��]z�=S�S�5L�Q�̙ca��\�n�.�s�Kr�r��}�e�ȇN�L����)��Wt���W*��88�Ͳ@3#Y�9(��Æ,�9�YbR1w��P�����A\#m#�$�9�w=�`}[�4��jkj2'�*$� :����V�ش��D�|���]��Dư5,�w�#�,����TZT8%̹q���[x^p�q%F^���׏V���Z��V���g�p2|�1�$�#�{���4J�B������tӍ�a���lb�N�e�C�w4�E�NZY�7�1s='*�Au���߀p���-ւ"�̡v`�,\4`ĵ��$�b� ��@��U6�b��޻nTV��|^�.2i��f��9.1/��9��h7iZkz�o�{4"�E�o�^U�ܜ���<�W4�Y�Ei���/�4�|r���((4�%`����`�Vq���0�_O�-�o�
��+P]�/�r�f괥q/�#!�	�M��E�ZsQ����z9}�a���� ��A`y.��Du�m�CF�����eC�;^I�\���A�n6/��SF���tua%f��#�I��9����a[��u��=
�x����>�꭯N��oO�����k�"�7��z�A 0���`k��֣��T��X�1;cB3���k^�N�	6��D�{�?$�G(L�_i��8^�YN5��EK[�ӫ��19���m�B J,�ֆ	��A���!��߀�y:��M�}�j�I&V�@u��"D@�@���{�3�j�����]p���ݽ�s�"K%'��)dsG��ĆZk��?῕�㫱�9���:E����Pl#�{�V�W�<��������H��E��vD}>a�[i��O��`g��}	��B�c;�|��,e���\OLMY�e��;J��!�.?t�������V��Mc�a���#�/K9*�.$x�w���R�!5_׾� �m����̧똷fN�����m���zDa�ux�/LfI������>��k5apu�󒄺z^%��.b�(��xi�Z���)H�7����h/	H�ɖM�D#��g[^�&�����[��5�G���S� �ق�^�P�T2Q��MĻ���k�&�8`��S��<��ZA����:Np�BU�/����{�YCK�}�?
�<�� ���_�g��S(n���d�sB^���F�S�g'oP9"j����Ơ������T��YoWj�F̹E�bۯ���#g�K׹Fh8�J\��n.�sI3AuTk8��q 1��"j�1@�:S�Ä@ݚl����"ث��$pņ>�[%m�׺��
�M���S�7�ç�R]��#�׵
���}�e��$ނiTS�D@�oH9��%��(@ٷ� O`5��gr����:?��K� M�X؁L��qv�zu���U��tH�*�Y���b}�R4�4*�*Z���[�~��kv�i�������i�����W]�����J��O�	?���+����
�*X���r���4���r��i�w?�n���n�fp	��Q�BM���]�!1�e<5힐���0d^K�⁕},����f��eB,W�I��_��&�#���$���kw��X"{ g��7�/(Mj>t혗�@h *� �,� XaVxb�7_���k�^�+�`aV�D0�U����<<MyPl5������<��_�3��0'�� �2� � #�d�,�`����;H�m�/�[x���9�&��B�����8D�.t.L�}Np=��#�~�r���k������H��:�E�[����\~N� q�,)��辸�ˇ����eȤ8���SL,-%��l�
�<�u>�R�cJ�|��=:������~UV�'1�m�0m�Q���a��i�'U(eR��0��x�JMG<>D�GT�>�F���h��v��y9��~��C���Nv�胝L�,��1���}��䣸K��ۜ�i:�K� ��o�)�- ��\?BwR��4C #��c8Y8��ڝ<龆@cө1ә7b�M��XR���J��e6r怺d
5��n`�XJ�P�H'�T���y�&��`�N��B�.�g��	�X:o��G�M�hA5���5�#��� i0O!i��T�v������,�z!�O���~�ͻ� �D!����ϞY wy=u88����@�⠭�s�M񃈦L"�#_�U@��a4�Ի7����d)��AI�{`��H{�6���[���`,�����@Y�<�ч��Gz�π_=��՝�+�BqXFc]���_�l+�2?Yr��	�Ny��C�����V��͙SJ��]z$�z�p+���W��Ik�Z��q��'��t�����O�{�GK��Nk
ކ�V�"T��F!t�� (��Kq`��Q	�+��ͱ�i<�w�� /Dg��%����+(ږ�X��F����e�}��1_t�ٿd��S�2��i *�,����:]��s�0-�O�fFE�8~�X̤_ٱ���M���
�[*n�js$��{}�V?���'C�W�|��萠�Bwt',��珞)��F��.l���7M�[�d�CG��)�k C��tҀ��������݄����D�>�
ޡjj}of�4^�2}hZjB$&��i�'����܋�E
};=�j�mo@h���$�tℚJ����5R,ǲ�x&�"\{���Y�ZR�����+4U��RqxøSS;���$�2�V����3���eQ�ف��c�5ݵ�pYJo�<Y����8�VL�����#���y�މ��}%m��UC��񩑌�eX�]���~���7���Cd���=��e�C��]J���R�疻˻3\>�79���u�v�P�&�ڮ�f�2�J�g�-l7��B[�B��FYx�L���v��h���Nf�7$'��^)杇�O�d����6�v�C��D~��?I� N���Ns���c��$@��~�E�"�I��^�K�=��Vi�6 &?}N̵� P�ٙ�v8���!�Z�K*�*�Mmz����Y3���?���o���|�Y�������,;��XJB�֑��#�1�Z�.D^���wP�-���G(z� `T9ѡ*�r��dSSG��(\ ��#V�J0�Gy8
.�Ķ�mbƊ��>:zj{?r�ԥ,^:���+F���\H������#���	Yc�)�!# ��\^\C
�-��K�Y�Ryk֒�6�̐��1�υc�9�n�ؤo�K���O�w��?Sߺ�{̉�`eP��+}z���̾��ٰ�6����U�����@99���{I&y�(��s���f��5
��&���_㈠=DϤ//��8�PX6�^~��hE89�����Q��v�m��J�2�b�a��Dް�,��}��l�7�NyD꫿�$@��L���k6}��Ve�pXr��jT�eC~= $�o9.��U� �D�
~I�y��H6��j�Yͪ�6E�)3�&����s�gI��J�5�GY^|6m)О��zW�nFf���[�檛�Y�����W	�:.5�P�k7��Hd U��I��;v>��?�	j���=�/�N�+y��:�Ƃ%����C��Yk����9P"�{(3Np���[�W��tEsL�����V9���Tb���ivG}�7h����!��6��j[�>[�!y����+����|�p#> �\A��N#�OfZ�O-ʲN�/R&��M@'����M:_+�.��x_���4����b�Nhџ�+�R5�t��P	��Wβa�WW�l)M�p���DƋ9ݛ�(:ǝ6�!�i��Zv{�����t��
X�۸��2{�`��Bf#��Y_��}�Å+�׶��3@ϙC���8�$?�p��l�_"S�l��3Z���u���U�]��4�f�s��ce����6��^��*�H]�^�$Ӈ�S�n������y����vou;닡���QM�>���Ɵ=ߥ�R��e���0�,Ǜ�BI�A��21����x��������%�͖*�,o���c�po��ߓ��J����f�]h/��+�\�g��n��
��rA�*EB�+b$�(�Ԉy;�%��O�,�������l�`�90$)i�L)]���O�R�K>�W�F�(�g0T9iʁ�F�S��H.zo�u����]����}	s�lS�g����ȡ�z���r�2�_�p��g������w�-�@;����|SqwPӈI+��bm��T^�<�%z�A����jJ��O�Cs��CI���G������� �����ݙ{،Us���_	Y��(�J������#���<�dg`}H�}
�	q�g�Լ��7b5��v_���J)*]{ Q"o�}^5�)�*�g}� ����V0���ص��>�n�@ͱ5��\lkuw�~k1�"A����_�ȑ�9��vM�׃�VIVq�C�7�I��ci�H[����/NB�m�Q_�sr���r�7��j�i�%wM�A��A�dc��z2v�B���e���9��|_��Pp;3x۲�����d/)��
���Wپ�h|y��W�]�OS�F�7�Nv�yj�1E���.��ow�8a� ��d|���,.7�m�ܪp���@P}�:e�¦�&Lt�-���]]�/u��q��_���B[��q7uH��9�X�;m�ӎq�XFAH�i�3ǽ�R6)�ب��6X����S�iζpnsq������`̎a�m�Ge�W��l4���~~�m1ݏuF��D^)K�w`���;v�Z4�r-��K�L����wϧ�O�l��M"��kY,/|�;_�ʧ��j���w��*���ǮE�\3���]$h���(�	���RxB8��EM��N�T@��j�m���ofd��c,A�C�Y)=��ʱC��O��9����̓?��x�F�����6g��44�h��ȵ���`7_|V�G�J����	p�}��sǸ���f|��dE�*���P,�ݧy	<�Z�wt���;6f��J�A�mU�/P0��HG�oj%k�Ƌ�-;9�Mt�on���5��4T9E��#�o�2���>�[V(�"��P���Q�H-+	.�*�(DF/nV�4�iQ�=c:(l8���6
��nLV�)�6��@`E�<|�OG<��g#������
���q�n�7�>#��vF3���߅o����T5c:�D��'>��v~l��'3�mɸ�t��*.�H�37s�6C��w���7��H�d�h�f�"/!�5u���{������QL�NG�z��M
_&7{��a@Oa�1�8u5�7A_��0/�������kWX#����#��(��"�>��pk�m���
�U>C�Xu�.���0��x��}s����֑�ǝE�>�	l����[�uC#
,�U��ki�J۹ψ��t��x�
l!$��l��<�J1��F���_>0���b�������XV�[h+���"��x�ɴ�;��U��S?Ȅn˧��i�>�!�E��|����GZkF[�����]��ʼ����#�T�?cc��_��������M�P�u1!Ü�?"�@�1�i1�t[��N��?�o4�G1sgo�ks�V/�k<� :�jt�`#_�����C nX� N
����C%����[��7 �Cy���z���KRm�w^v��ާ9���e�,g�JP�o R](��,�jT�v�LQ�,�oZ��ڇ)��C���K(���c���5M�����(��������}�y��^�U�8�:f�o��@cm;1�o\'1ԟz�M� [pxXC�z��e�z숔&�znXw�~��ho@�K׹>m�����-x��1��o�yf�\GK�]ƃ@��#^MZ�����?���IJJ߁;��b7
�Q��ݢR\��H�LFA-���<� �9��Gf^��F� :�X���((�h�	���n��dl��/��Q���O:2�X.�Hb����-%2�Ҙ��Y=����qr�+w�έY����U��j�'��( m] ����a��{���|}S'yE�:X�L��]3��O+-�^�������,��([�DI�j��xsC�i�M7�6m�
'�u��$��7�c� �h�խu"�M����M��?�����n�7�����F�`�Y�#�3$�.��k�.�oJ���k~���d��{i񱪞r	�P!8��<,����^bh��(;��/��'������3�����}73��.X�Ԛ��xRcgE��\p8�ʻ��8+�ݢ1�	���~]�]��$��p`D(s���2��W�����`���	aB��[]KRG���xQ+g?
*���M	��}F:kAEVT��bư�5�� �+/Tˮ�R�4/�F��}T�H��8w2��Ah��Ih���箮"�)�~�Wi�"[_~�溎yݝE������x%��Z�tM��>\�/A;!.�����
/ڔ=��0<�Z��X��-c*Ưb�`���^W}��������Y�p.��2T�
0��e����D6.�Rzčv��T�]i)�7������AV6�} �S� �2�OJ|g-4�G�|4\�Q�[ѡ�E���bë�Z��	��w��㖷�3Kn��W��>d��tE�HᵂWm5��տ�xE݇�*n^�����EKnP���>��y@�p���.:�biP��>��u���
�^m��#�~@�T��B��Ym���M+S@<Qh2�$�&վr,��62�@i�vU�[����!t��b��#���V!v�A���(������~^ ��A�vF�7VJ�fڪLf�"$�O�}@8f�(�&�m\��˿��c�G�x��qo*Q�3cQ�9��cKN�T��8���oE�*��۞��ӍCӀ����<ҝ�2,��ʶT���@x���(��H�e���?=�2k��q�>�.�Q(��Yp	g���j32LP��^C�p��q7�g���ZU��զJq|����A�r�x��a�OԹ���8�$Ъ{hĠi�/��z�����g\�=Tq�_殁�a�A�Y�Jح��ʔ"p�k����M�r���	p�1��	��QEs=W��'�,�7��t�̝�5,&9gt��3}��A=�V�tC�tטߝ�Ԛ}�	{n�ޜ�`�T�H�\�?�2��/F����9�G����V�;H�DP)�n)#�61�3(f{_�f�c{p9R����L�T��V� �bߗ��ͳ8��7�����J���ٶ[�b�e� �4r�6Ի�j��M`�0���Dq�fכ�a0����1@c@d�is�o	Ζ�~� ~|��
1E���$:Ư,�����b�=%��G X�i0(������Ո�8CY^<@�����#eȨ�4����q&'پr���=�ۚR���L��RS�JTEÁ+�<�z� ��s��."����j�R��"G6~1�շT�$�Gp�ۑ��LCaKkJ�xb�_}�:Cᙩ�cA��B��-��u��=-Uz/�3��3��fTBEwk,��25�6��:�����S,�h-M�f9�١y��:��G���#�u�f�-�&I��;��ūV�T���8�C�u�ߝ��IHH؄[%�A}C��{�� �|=p4�{sxs����ЩL���_��,p8óu�M��I�֨ae�.�K�Z&�|F>��9&Ź���R�C�񫡩{=�F��yT}����U�?���� =��}�1h�^��}���L���1��yBu�Ml|ú��Y�8KrXP�:��E�#��r��z� GY���(��m��K���T��8��S$�r?��g��G��1� �X�~��,3���4v}Ѩܵ��L�s�0Ljy�즖�(sJ �d�zT-����4������$K<fl�������Ҏ@�œ,��B��wb(���s)8&����I�埝w�ż�G�J��� ,��>9���ΝmM=M�Ir��8������6�6,6�vF���Εc63�����޲9�YF�8�� Q�Ҫ�;Ҟ�x����� ����������	٘e
*<ߨQ=P�bBU�޿"�Y��
�Tֳܤ�Xk�+a"j䱺�H��S�]W�5}u.��JzO�o��W�צ�I!+�O>ʫ����9����&����~�G�`�
�3<�JF�d ����ie~j���&�pD������+5Rsl�G�Ϭ]�Co�/��8Ssf2驰�s��(ƥ���<��������ʈ7�"Y �}@�sg���dY���5���\--q�(�>ܨt�X�S7t��+:�x.�X�[����i����J�4�A��
��y�%�??]��޲	�Y����B/��S|���_Q$��ޔ2�=���V��t]��s�'ˤ��X�Mk�I%;诘TI�H#;�-BЮC�$�K�5�F:����f��a�}�K,��U�vh
�&� ����edGT
Fw8���sC�9R�,�X�c�K�=o�`2|J�#a����*����g����l���Jɀ۸ٳ��p��½	�c=/����1
���"��U�U�JM�w����sx��<yFѳ�0�$s�&�F��1��8�Κwn�U����%�5�QDD����,�^�Nmj���`o�L��?؝l{�ŕ��x�JR"1`���<{�*�E\�D�]c����k��ځ�M~O��>�"��*�e
m	�����)���:�6�8EͳT��Z�1��^fa��y)�_90�p�a��:�#��WC��(F��?ԯ�"t},6q��j|��%�8�L�▰tϴ�SI!�{o�P/!�N�+��s���m? �3��!���JTG<�q/�f�˼Ͽ���:y�$��=>|��EA
meUE��Z��7%�U�aE�(��]t�)1!��!PWc?�T�f�|}P�q'��`�'�(Ȝ�g I�;%����ʈ`���P^"9oMm���Ua.]?�4K�w���.|Eẅ�u�C��¦�ŗ"���ч�A����
��Y�$l&�Ĳ�<�-H�������[������G4�XjY��K��^k@4-�l�����78�=�@p�,����_��N)��A���q���%��KJR��'��&��- Źdkϑ!��y�X!5�䌷TQ6����g���v-y8�*<���D)h|.`jf5+?�����A��YB���N�X�] ��&�#�k�,[����>�q��x/O>��X�#I�h�M�&*F^t;�e������E�Y��pR-Gpgkޕ_и��\�m#��oޅ��H���9�d
'��w�>E׉��ZP��F���Y��g�u's�&��~9��;�/�Q&�a,���F���T,r~��.LyY�cC��0G 
�)!��L��B ��/����yV�NޞM�x_��گu)�c���b@S�&�oLT��GuMG�:]׭�3+/U����G��^�YX̒�fo���ql&�:G�?�#��EGH�2JIY������'���L[Q5���)�~~2���i0B>p�et�3��5f�m�̃[,M�7��i��AeX��Bk< �!3��*و��e�Pm<���s	'�>�;����P$w�"���5����75,.��^˝4�K!Z؁V�XΞ2t��3>���Wa�d�a:~\��PQ���� �D�e
f.�Se����r8��=o-�^[|�׍��Ԕ�/��/�50K���A���!F��X@E�!"���q��	kos�
����]��kb����-_�2<�����}6'������0eݝ���"=���jEy�`��d��yK�@��(zQ�.�������P��j?$��v�t�ݧ�Q/�h�A�Ii������:�9��Ksg �����
X_���f���&���O����z�^�� k��� q~U�Ģ��C��qF�W�4�����4	�<%6@�f��_u*�����Z��&$c���dh�Ps�p�GO��(�	D׌FsǪtE+0�kg_�hp��!��+�
E#u(��ʱXh_��l~m�&_�8��l$���8��p㢙�O*��v��-�;��K�^4��M�8��HQ$�N#ƅ��v�[\
�����$H�h���?*��M�/�6|�g���E���c�w�3�\6�a���6&�l8^k�\�q7#l��t������Q��>I����>��{ �3���i$|��4�|)m��t�F6�4��(�M�us���b�c����>���y˨�1��\�P�y��a /�l��%dK� ��)Z
"B��G��H�v���X�K
eǎ @�K��j����ǂ/�>[C�'���9L8�3	�����5X(�{���[4�,���GB�Cڈ��E�K�3Ƀ��\���\�r����!�(� ������7K�|�f�ܖ0�О�<"�VّYu炍V����vX���K�&@��-{3lVI� ����Sc��G>����-"��P�������҇�
��G��@y�x�]�@tD}%�B��n��gS�Ol�,�_�@���T���<p9j�w`Fw\ZA����FJ�RHe�]����]c|O�3ѯ2AS��9ᘗe��Ͳ)pd8 z*�oK�mw�����#��-����n�+����(9W=�i��$�7q����E�ګM�\��w�u����
��cߦDy��q8���j���G�EM����n���5LR�	B�t��M"�����9}*j@#��ĳ^髊��v��x�ٗ��s+�ٟ�2�,x��S1�����ˇ�ì��%a����\�� ��ā&�ѣVj�^z�I�{H�	#�(H��d:����gf�F��%�(}�����$��&�j�̺����_R��XH\�>]�d�!���6]a
� ��r>��3G`�;[��;3��<?�����SVs=��O���u����C�t�ޓ9�������E��pO�^6Z��Hև�׶�@�zd��k�7ם�\�;�L�(�.�7��و�E4���,׷e����>�`]2��O���{�H���X���R��� �[C�N{��R�
�T�S�7>j|������R�a����h��a�݋�лN�_� ����(n�K��n1��օ�rVD�E��Ӆچ��gB~wϨ-3��k�x�h���#�#�]�^�b�Ӧ�ȝ��0���1�ZG֕p$�n���?�z)X{o�{�Q����u;z��uV��n��a+4v�����O!x"U������?�9����TG�y^�C�R�C��N��
�w�_����h��i�W᜹#V����GmT~���[*�D�JM����<	[��\.=�x"Z��i����^��H���5o0��=�a�I~H1�#��{�5����;�kY �M��
�d.��S�u�~M�Ԇa�޾Ak�R��Ԏ�ַ�C���֐��>&šs~��5Q'B�C}����}E���w�C|l���z<��{"gv�O=��ǩ;*�M�"�s�K��]�q:PZ�
Ï���w���ۉ���=/��CS���}#n���l x?|C)�{��5�C`�
�5"�)Y/ى�k��L�&Z�#O���	D?�Dw;o��Q�S)�n@��3�`���ؒ��7ۘ8�����+/�+�"���M�8���L�zx�ѓa�����L���(+�e[#]E��M�Pjt�T�x5{<`nz|�]#v[E������qW���u N��O����m(2e���\[3��N�JQ$Y�����^~��@����>`�WŪ1|k���1��%�s����-"F&�C>�h�4� ��肁�_=z����GGW���'I����'����.�� ���^y43����@�O���0�DRK��P�`�R��/���x�<)�d�ʻo��Ԍ0�g�ɾ��{7����j}�G�#Ĩm�aN����Ӗc�9J4��<�zц��:º�*�[4W���(T+.@����nZl�۶=C� iq!m��o3��}s$����R:�`~�q�m��A:d��L}^zUh3M���nj-j��l�_�Jܔ�>�|AsGkl��|1��Ǌޫ��H��]e���~�o���=,����|"�*c|w@˒��w\v��f|����9���؂��b�6�4�>5�~c�V�R~����&��]NX~�B�\��{5�9�R������z��F`:kY���럐����۹�)�᠀��ݝO�%��Q:�=7���m!��aB�f9T������	;BҚV�l��^!Y��fo ���x�h��ҿ��2هB
ЎĞ�_)=:̠e������z���u\S����ܗz�g&.0�'5C߶�����uDxcN�ԥ�������d�_,\yl5ؾ�4�`���2J����<���pp9�1Y��E�x|��{���0uD_�������l�J�I��0�AT�PDo��:+	��b�d��\zD�Q{7�^��l8��Z5��)��=�o�;u+�'���1��7��ծ��4Iݦ[��W�|��`�K�0�
��0�7Sk��]���9�;v���N��\I��ҳ�7�8��b��g�� M=��
���K7tƥ�����a�������<� ,TA�ph\�[ɧ�2#fң'���w��_�ctu��l��9C��K���[B� ��	M��-j�da�P�q��%K�A�R�n����<�
s~���߄K�+�=#X��az����C�?@�ҎF�1&b��jy0ͯ���&�JQOk$�� �N�����|��b�(�Bo�Dz�A�&Y�#m��F2� ���Aw�;��z�mO�����_�:��,Dse�Z�I�����_Ac�
��_�U�����	k0�-d(�EM�|V���'0V3�;U�8ÑG`���|�=RL8��U�(zRV$�X�8ؙ{Qs�0�h������('�Q'�Qg����jIQ�~B@Hin��C6�Bh&d�GUTD��.7s��\����PM�]�p���p
v$�_�A����s-_i�_qǧ����ڮu� �T\�G�Ე�����ˠ׬�+ѻ�T�)���>�	ņ�12��s��,#� ���";�	�osb���
�tvo8K�x���l��/'cc^��3f�	ePb�\�Z�q��(��`�=E���ƝC�K@B�&�G�h�������tl��V�#�o%F�$����?�P�e�la��6gK�a��Wpe�1#��7�1���\m/����a�O��<n(�z����z ��n�wSܰK���^��Lە�F.:�B��W)�2���cW����������8�Јf��bhO]�gX���y�ӭu_g��!��J1�i2 ����?��@�]/i�l�F���ku=G�Ԇee�c�������.�Q��w����J�o�C�������
��8\����'v���}�]x����ڴ�m�����<�����b�TZ���Ɣ<#�h�����὘��Uק����E3�x���4�%{5��X9b��Z�<?��?�Kc<sQ*]�D����V���Y�����{�{r�ۦ��Ǘ��f05A�xp���8R�9F˯�v�����ᬸ����m�g1B�eJ�A��j~��[A	��ϟ���$�������7����>�*��H� w�hb?�0���[nrav���vK�����Pw�W�T\��P�����
�h�T���ʽF3'���K��jt��6���g ���yަ1C��|����8m{%�?X��WPp��K���s�l��x7�48�'�L�
��fY�k!��q��7Jy��/\k�%'�=�I�ɴ�MT}1��8i6�c��yR��bv�A��!v5f��b��w���!#����e翦b�)�xO�a�닝:�yL �#%��E�3���2zF�#K�4�#b�9��t%ɕ��]�mK�ԫ9�l�Ǟ�I-���%r*ƌ�GՠT��h�v�V��բk�6��ܝI��y�� ����]�r�U$�����b�IAu�
�,~���3�j;(z�;�H���x���%F�n��<G8jU�k�˽�:�ů@Gsq�$��y��4�\Eh7�ѝ�\,�'�ɳk���9H�lU|�\���$�x�綛r���'�K놴�bƓ)O����sq�zec�W�%�IH:)�w�Ä�V�V]�%�j�#�t3��V~�뉗��7;����E�j�i�������ɸ� ��݌�մ߉��%��� @��¹�sj�^"��W�Kl
��L�:e��%z��Q�#�Y��m<�p��mU�dS4�q8x6�`�/ߒjz�сϛ�d�+�T^E��=�T֒~�����ϗ�rX��Ub!�r��1ʮ��N3�P<q���t��>IzBR��kWt�m��>�hA��\�DZ�1l�N�^D<��Z��C4!��^�9���[���,GѴ��GV�C'ާ9[U]f"�ˣ�-��� �+�թ0�;v�t���!-8���|��P>�q���n�W��w����(�����(vn�N���z,܎gaV���is�#H�2u���:���$E���:1Տ����f/icPi�Pv�0�z'�E=�!sYǶ�H�4"������"����/�QD���P�`��1���O�o�]�R@��������r~�<3����G�aj�wx��V�@�1po�}G� ��|�(7饠������*pm{2���X0�ML���[��p����-$v�>������#��TZ�A�����Mk�v�p��a�Ӈ%��.�jF@��^.�o��͍ąy���}���T7��C4��������r֓��0���LU`wE��t/�i>[���T`�D�C�-�|���T�պC�p�F��L�����6����At��k�S85��,jQQ���Ұ����) $��	�%٨]t}S��Du.Nb׳?�Ѭ��!�/�k�o����K���J�Pi��Q��t<���<�	�����:sڥ��2�y��5_��o�9�n�KJ.v�W`��&=�_;���2�Ϗ���&�pW`J38��`{0�nZߣ�%q)�U�@����1_{��(�o�$�v�RE����K�Ye��o:�_����SF}oS�)����xo""���hz�ٓ�(��v��'	�Ѵ J�5�Z�>&��x����@^?"	�p4�F�[�8�S��,R+""�Ҏ�ӭ�]ި[�oMS���*7-&mS�x�k�gS�&��Q���u�2���L�WFl���'@c`����JU���c�#}h��G%�3@�U梒���Q<͝w�G+_�9z@J:5���H�P �ўRf�6X����vډ�,�P&��#���Ox�J��uto�)ι�y�
��sL�)S��ʆ�`��$!��I6q;b+��83gl�4�^���-ViK2c{|ג\��|�ǲ����u@�*=�>���U����r{%�[��MVj����T�݈m��u"����s-�}^Ā]u.9Ĳ.�{�6;�y �lc���H�"J��9Y�5Lfg�ʈ��#�Zb)�ɜ!��qɡ���Ƴ�pŘP�s�|͐N�j��,�gA},�S~'l}j��s9H� (��N����s���:�v�`P9[%��Z�x��(?���H�2�E��M������n�~/����	�J���|��4��>A���@����#�C�S�h�ڝt��-�
�u��|��I�S����
 j�j����`&=��>��]J��G�#�XV�H��>b(C��������DG�l�&j	f���UJ>d=q%꽽h<~Q�v%��Q�ј9��Ok����_�tHu�&�������1�Wq����M+(�ZW ��h�a�|���v?������	��Æ�j�xyE<�Ȗ��O�Ǧy��%�a�@Ny-ݻWRm��gRpҀD�fWVT�]p����F��p��#�c��(��w�ۻR[3�t��1�Щm�쾓U�k�P��I�K�e��t�`=d�f��4:�����Zfe����!�ʼ��XT�,��ڄ)�����.=�Vda�1�
w!)���&�Ƌ'�,ɵ�x�<#��Q����u�	w h__�:����sҡ�M�R�]��� �������*��%��
���ͻF�\�F�^c�C#����k�J"d_�C�� �18��!��Ks5*�;8�-����m��>9�uR*m8�!�:6�4�,�ֱ@T��鶤�8��x���rO�_�Q���~�u�5ޙ����"�>���<�Fkщ�ϰ����+��*�h���%>����� �w�X�aO��=a���k?4@�cVk�="m�f�%���pSSK��߫�u��;z���810�_����z�qp`�I
{���3��R�
ap��(���sZ��n�p�2b[�.7q��ђ
�n�iV &�����TD�<�q?��X�p�a�m�W�"�|��a�ܢ�+�lA5�yƎ��ȃ��T]��)j8Μ�;��f�����2~3��U�$s�)��n��
�`�;��d:,{ �:�-����jk�?�J|ȆR�ⱸU$�B���������_*�]�s��_��j�H��=���	.��V$x��wV�0�O��H_��W���?���>�dS*���EZ3$�$�\����F�d���^�J�O���Ք^��4;��VT�����h��
ŏ���Ns�}�����ɶ�%���u*�;xy��B��i��qqYے���M�!3�6��`cm���-WG(7��dAo8�:_Y"�uJ��K=c�b�?n���Y�7҂�`'�}X�^ǌ�XŹdh�e�ܨ�Gi�_�<�ȾmXci!�`�a`��B1����5r��{V��",�Q��6��S�U���~X.�O�CU��X�i�z[.�q���$\���Q��e�92�M��t�W#��ܐ�������p�Ǐ�ߧn?}��&�q��k�/fN�G�ͼ#{��uY]������C�W%����dq��k�R����r��'�6�Nح�����r�5ܺ5����[|��q��������ߗy�i|�v����A���G��]9������nx{�"[:ۺ���;Z@��L�Ta�S����_+BU�Ӂ�x9_er�(e�_��l�0�"ѴY]K[.�����Z �aQ�HF�Q^��2A�2~�:�� gh|` 0E�O��ʈ�r,�ؒ��݊�_�Q���p���H�>ͩ�=�-+��K��c��RD�0��>�v9-[��EK.g���Y.�����Z��i�O!�A�j�����A�o&���b��5��n��]�@�a��<���.��qP~a�{K�qįV�F��Ż����M�;���q�EuN�8PZ�Y3�`}%{���pd�O~n�{^��o�t���T� &�Qi�F�P,_B�~	��hs�'�2�M�7w�
���x��0�(Xfꋋ�>M�� G��������X�����K6(�e�()/���$��J�$���� ~��&~Y?�����E�/�FȰ�T
��g��ڙ���~L��o�$	2�饸��e�]�L+����� -A�0Ϭqր�ix�>��ͪ�N=|�xF\jx^�S�Q�`wD|����E�p-���1U6��׏��j��;?�3�[ʌ�]�ц�%��Z����6"[�\5>�W��yx�I=P*����v|�6r�����x�k[!�8�`Y�����T�it�1��=�\b��5��w���zv��z�
l]�"2�(1v��j���ln-P�_R�&��@��y�������m6�}h�B#��|�/ O��>5(���p�F�]�޲ɋ��A�����ţ��OEHx�7a�t������*JH�<SҹZ[�a��.`M�Q.%J}�b�� ��j�4���O���).%c+�k�V׊�^a }�>�t���ɷy��߅ٯPe�ɗ# ��ӿ��2���G>Gھ;��s�{0�d��9��,�j �Qq6�N�1�{���#��v�D�lƃ[0%�Ju��Cq�Л�O�S������"0�����_��D]��$]�6 ����>Xl`׻�	S�)ۖ��tԷ��:[�WZB�}b;
���z����d�uo�[���)�x����w#��V�,��.N��r�`u���8f�r� ��3m���^�)}�y���J�9J��dN�� ܨ� ����ʽ�Ns��H*�$F����y��>k�鵘r��"�.�_�R��T�	k��L�@<��FA:������q˶}K���8��$��'��0#�:���W�$|m�]�:�ΊX}!C�n;
N8}�i�]���uyTR��. �a]K�S3�^�
f(b�*�����mQ�G�c?
���y]�����zr13�`K�ݠ��|�9=����6��Kԝy�u��Ԡ��CU����MW�W}�+�7�ll}���q 1|G���4e{����+qc��̅�ߕ��F=W�
�vkx������������A&xNiD>A���C;�0�1A��K��Uo2d���������ק�G��B�U#��(#٫͇c yG�b��[�W��P'lU����sv��o��*���̥�ER�T��S$�؇ċ�W�Ѭ<St6+��BhWTr�2��&�	��l1C�}�_ř2K�������: �"�]�v���w]%�ꠕʮ$��u��E$q�e���ÙxI���v�E�Kj���D.��Gt�+�>�D�Ϗz�ٔN��{�lCq4��o���c3�;�3"yh佾�#&�0j�[�%E�u8lWqf^�e�;������ ��x��H��*N2�}���/33���#�\��)�3N�V�%D �n���ء.N|�$���ܞ&�9a��*-�q�/�����=��e�`R,˃\c��,��+�h|��ס�Ӝ�<w	��I����g�/#��2��+�f%[����
�ɗ�����q0UD �&�M���/bת��w����T%�[�,�J�֨�� Z��T�]��ߒxo�)vI*�DX�������m6feo,	������iYĲ_2�}$��wK�.�J��b�+׀W0ѪF��5dXъĵ������29�X�c`~X�he}�o;��C`��4����r�\����G��ͤ�[L����C�����k#%��k�	JD�e[����t`�x�Bw2����&C�MD�����~�H}]�^��A������ꘌ�u��S=�pez]�A�.<��l���?�m�/(<*��Z�' l�ʚ��d�P`R	�懳�݂��E$�a���P�_+'� ���괷)��g��u��\���Ν�����ܷ4�ݱ�G?�C���{t!	�k�_�^��9+A5ۚ�����w]�0Y��K��߃rKMX3�h�f�9�2f��?��)�}���y�i��6Q�S�X�"�<�6V+�����qW^�3�t���&�w^ݨ��H*(�Ÿ���#��]p@��7�Z���bi��s�������X���z��݄�;��ϟ���V?I+��ݺC�d`w���k�mT
�����k?}�ޥ,B�����Gyl��qJ_�X[����p�M=հ�7=n�|���͹�O'} �7���B)f��k�����k;2t���W���^��Ŕz��8�(yǗ"��@�sXs�TsS8���(��a�Ȃu?Ƿ�`��֐{p$t��wY��q���n�Z����U�^.B ,�!j��bc�D���)�1{��;�x��=ߓ����MT�n��6�b����M�"�;j� M�j1�]8�
����){�������&�?�BZ��
F�A�8�	.݃Hy�'�vM�$o{��:�����om�6�4�����t)��Z#{w���Fm�<�t��ڝ�%�*}���	�^s�yw������t��Mԙ���h�=sh����.;���g�"����UPw ��Ϟ|�'6�4q y�z�c�k�\��I�{�2�U���s��I
Ѐ��b���}��k*��u亐��(�o� G�n&Bs Q^g��.���.T�l=}&�}~Ó��� �X�a�M�!��=��
��B\Ic�%��{a%*�!<.��=�ɢM�L��o�Xye�z΃���6�3]�8פ^T5��VǤ�ʡ�NG����k��L�C ������,�_�%� ��)�}��
�r1����0�~K�x���d�����ߦ��4�̭�YS��i�ݨy���Ȉ��w(y��t�������	���{mm�؍�#M���P^�_��'A��00�}C�Hi򣕐�m�'�����?#@��k��1��a��r⛃P/6�7��N�����Q�3=��K��73���"U~��B�@GYe�Y���Vzz��'�( /�-,>�*xe$�C�.!�,n;���vw��i���
������0�d���s9�w�i��2��ϲ��$:���1X�������:2o���|�_��f&�?���5?�ǫ���[������E0�����X�I,A�V:��=E��9m�  ��f`��fe�ahh�t|c�����o";�NR���[/���,:�>�H���sg,�|)C0=5N�+;h#�#�7Kɝ�KX�����!��Q���u"���%)�ZU�f�W�9�SKed�I/��t3��U5�m;p�����z������Х�
�W�E���{8YN��I�c.�K�-���{i\L����$p箢aI���\�W��Q/�ؚ����o�?	��f.��ʖU%d�c_�l�	lҔa"]F+�6�[�3JcSM��J��'�ro��b����qѬ���o�p��;�7"ib��񻋏�2}D����8iӼ�Y@�FO1��	Q�Z�J��N^z��7��U2��L� �K�x;쓻��F�/���ݟ4�!�����)Z�Q�����)C����*^�`
�|���-|���ͧ��q�dqVCq����COϼ;�����̈́�����i�3��,�7���S��~��9B��`?�(}9����~��L`��U�Ŕ-ҥlI�<V������7L�g���]�B�$"�=�#�H���_�pn���[Z�5�a��Kl�[EN�������ڲ�k���G������]�e�Z�DϘZw"��	`%�n�?ȣ֡�C۩c�H�Td;5��WE8G5ˁk~����b�K�iT_���W�!(�Ȁ�e�{H���%>�Yn�PL�^|��Ldȭ�Բ����k	���}���M�xcs"�\:*�&�{�`�e�n�jnA�,�aX{�y�2��Ԯ~��5���O��#�%���K]���X��G�NChM�$��<)�����᪟}�D���)!�.Y��1==�TM# `�$�|�(;ޫ��>�r�-��B��IXV�`��Mߟk���� ���C�+�� 6������A���R�}����n���.G�&Al������굔&�������*�Gr�C��ƬT\��o�f�:D��������eL����MR,����b[�u�Ҋ/k �*G#��E���K̏W?�D�xԆ�y���h9sǅey���?V�0�8�����9A�CX���?Lד���[	YV��e�c9���b�}�}֊ј�c���&P�Q�V�4�P���(�Кz~� l�>Y"//hCIoh���&����Ř]Z��'~�Y���)��?�4ɳe��&��H�a K�sW��q���зq��Mg#Ά*�G���3��L� ���O;�� y�zk2�\S�+'��-����u�7�ʇv����ŕ.|�H"A��z���%����h�o��t���c��?\<�-���`�� In��(r��%.��# �
�[�Lj1�q>�H��,��97�8�h����U6�v:
�L�<bޑ���PxqG!��J9��ӒN��"t?Å��.-��͉'��S��^6��έx`5��3ќI���qM�B$�����	��G/��_gV�>��aK��poK�2O��"�zc��s7&�*�Sȯ�:��ҏk� �=��!L��H����xU��r��O\'�7�sJdj QnA�i%�R��V��8DIN����{��ɒ���YF��;�hOD�\������
�-.֧���lKq��2�6a��<(i�F_�x��pF�� �r>���O�[���	Ȇ��K#^>��OZp��[�����I�� Ȃ���b�D��)0Z�Ao��:�h�ASo�CE�!���iJy\��\����]S˲��C� <_�^h�WQ���8���wv���Wus@�)cS1���%N�i;�0�� LW�B�io�{�[�AG��S�6n��Nt�t�����9_Iʾ�����Õ��ePIyj��R!�����OZޝ�"��Mx�^B����K�V<�����ÁJ����J<�ؐ��⇂R ;�N>��`�E�A�YE{2�zU#h���VVp�r��`'D��'G����)�7m��EA����L2�ƭ�W��"y�I	p�Ok⁵����qN*v�Z�6�a�P�17����U�^o(�(�U��n�l����8w�V�9n!�)Bc�1��Yd�3�)�k�!G	G��~8 Mdq؞F�c#��S����T��y &�#X� �H瞼����GY|��ج��I���H5�N]_�U(�*�x^?~�=�RU�4�&�h�W�X�K�=����O�2&H��ba�:������yתҠS�^^�!Ӑ�[ryF�Q�l�{>�ZJ�z��(ᵐ�
��k�	�gO�@��B$���y��Cec��
�&�ժ!Z���ןzutp��.5�}	� ��w��+���D�2�AH��7�|���1�����s�ܾ���_�5ە�c�ثa�&����$r�Fv�1��,�|�2 Zm�\�t�ya�|���+6���U�Lq ����P�B�N��>t�q|UG�J4΃	q�Ev�x�I��3�i���w@c�0�{���j�z��J�
>gv��|��j;]n�O�̓�o��<����υ,��U����)��5����%;�W�z1�^@L�!���fM���3�HS����5R�ϵw�k'>���^
�q�'���N���m{�.Z��E
dֺ� ��@��|�����[P ò�nC����W6���.�)Z|V^�Y&wS����'L�2+U��`7��f��ߕ���H|"k�3EuC��Z����ʚ�BEC��@�&�؝9��5P�N#��獲\WC$/�?}�Z��s+��v��� VrP�`s� �i�Z}5D<Z��j��й��W�qG�J�L��F�XߜU�H��g=��5vZ��G�3�qM1|�2��<�R�UU��z�	����7B!��BJ�(u��Ԧ�����N~��[B�ݦ����Z�$�*s؁ҍ�4hyz8��Y��R	y����Xp(���~�r:R_�,��u>�־�+Dnۜi����L�E9M�vx.���T�� Z��$�xe��m�A�VKU t��h	+ֈr��9���q�e۲�B�8�Zi��@��;`a�G- �d�Y����(���N=���>�Q��/zگ�(^������N�|�'P���5;c�FXu*�,	����=7���^Ta+���JRJ�@9OM���Ɍ��rDp+�M`ӫy�0]dĢ�Č-�W�;�,�A�_���������-�|��ȳ���z�\��t�0 ��pUV��Ա�M������Ջf�����N~�����X���n�ȇ�xJm�,(ʱ��Mj�riU"P��A�uVr��>��c���]
�Ź�CڨH{�F{�M#a�V%�H��zX��fʾ�� �����*�H�/��d�4������E񂖞ֳ�"/I�63�]�����G��A�}�,~�@7x�|����
՘���mͤ�زt�bVo��Hf"��Ѷ��d؏�i��_*]�}�m�D,���c�Nܫ։-��I���wti7!����mHt�řt�|T�1��"�hըm�Am���f}G	�M�r��Z�9j�z����ΧLѩ!<��-4y��i dc�pM��N&\o�G۸�����:DjK�pY�z bdfV��7:j���.�����4-�����o�X�)�����[��K����g���k�)�����P�s���CM[x�y�Q�����`ΉR�R��O�.�v�S,����U����9Ή{�� >Ylb ���"Jq\u���n�?�@?��F�:���~u�3U��̞��E 躧M���]K�E�/��������d��_{��j�,�<W��=��c�n�X}6�ϓ���gr	&I�b�/#����d��˄U7|�l?�y���S�7��D�*����k.�Xz9��06"�[��SN&]YV����Mɱ���9$Ǒǆ�M���w�T?����DW��_!E�F�εڮY��x��@)e�|�1���B���΂�}��vd�{���(���Dv
��\�g<6eY&����+���	Ea6�.���b���q%c�Xt�ʘ}���ۡg�i~O������[C^j��,cn��|rm�e���A��nL�(�@���!�)8>�qCr~ r���Y��E���+5}������u>������Zz�@6%D���>�Ws���ʹѨ�R��P�ǋ��.?ڟ�w3=���h����)�[0b2qe���*vY��	)j�c- ��T,�$h�{3�(�bC�+w��(c=�� �{;��E��F�\�i�q��˞�XؚX��#7uN���w�Cׅ�:�U��U
ñ���L��E�E`��e����}Ђ��~��_Tid�Rm䐐�����ӥ#�ϟ�כ�N!c�r��E��eD9�����p�@5k:S���6-�w`���Y��#�����?~�6U3��1_i�-e�<�F@IO"��v0H7��ѥ�,���sB4�8����D���P��F-��������9����,�Ja����������$��<�i%�2b��nKV�<�!kT���p�<!Z��7�י��T�J21ekL�i���O��L���Gpt���u��)�Ov	RE�*����1c�L�fh��#o�\��z .
�B��#��K���;� L�S�x8���s(Mɵ�!ZZK�Z�h�	8�'f��$� �x��$Gv�xȦ��p�fvh��>ݰ��	M�"�/�"�`;*:����jh"k���
FoHJj,�Q��&�`"�3Ӊ��c��\]��M:�q��  ��L�>�R����p���.�.(��4����Z�Ë>R
)���wiI�o�gLR��+.r/���l�1�/(Ǥ�}�w��t"fY�+��`���_+ȟ�����p�(>�_N��z8��:)'�k�����w��s�Z�)N�t10-A�]��Ѩ�B�g�S������'���eZ3�3�L/k�h"��u��B���-.������-�t!/���:ڝb��fi�#޽������Kh��Q����rOܬ_ˮ��������n.͞�&�Z�,dh{�G�+RV�x�>�!�w��(\}���&���3[;hf2��W�㹙�ʯ��vJw ø=��΅�K����2ߎ�Oe�L]IY�~�}0��j��B6�=�P����*c�A)�ַ�ngqèވ3���0��B!Q��6a�����zj��7�k�ou�26t��"�E'uP��TJƯƥ',��D��:Ћ1�+ۈl9?�̵A�nh��d���m��M�n��_>��a- �ŋ2��������f�@#7� D��[�p3��s^%e�Q���a5��5��,k�d}gi4 �W��`�qKr�d)Nq�%�t��� F{��B���g�ĸ�rFf�}=��I��޻��%/4b=�)���C���وgJ�����]ӨD8>3�oGl�u*����;��Gz�������`��x��K ��r�^�c��j�)�D.�v]�ȝ�82�&����2�"�Z�����OT�C�r��L l�> /&�uk�M�T��'
��\T�t\����ؖ�%˟Q;+��z2�˽��Wk�(e3?�����js���u"�U�1x����F��>��Q�s�]���Vd3�@����`fG��T�������FrZ~�}E�,��p��)grb|��&�a{u���D���?�Pt�N0Ȩɲ< 5��a]�~�}7p�b�_W�Մ �>�2Ϳ�\�y?�j�̲���B^��<	��]����j�U���!N;�k����`��jת*s�)����EmC�M$V�@���>�<���.�T�Js��R)�qkqƆԋ{�1�D�k�������8/�Q��j�;���:,���Dof�|����*X1%uS7�j���FMz�+;)9��r��<�|�v�qϓa�ֲ���Ex#w(��>;g,���ʆP��Ns�512�1X��ێ~,��חc�,������|'���녯��E𗶯��g�8��bH��q�4�S�E�TR����ў�铋0n=�8)�ࠤǛ��o�nN{���*�S�t�&��K,�%~��s��uk�]�~����=�©�GM��HF���.S5��(��Bnj�.�3�^��9 ��3�e�m��F:�]<��zd�tk�0'����l�={��#���Ig,x_X�~���W��Y���fJd��;~�&�菿s^.&Z�2��me݀���?��NR̩�O��(	����Q�b������K%�D !�:�pw��Z۲���@ٟ t�H;Rr*��W���^���\T@D(���'w��Hy��c����A�A��jbv	���(k�H�D��W\!)��4�q�ȏ��J��Ma�E8��ib'���OQfY��M���LR�JN@֦��_�󭧞�+����K`� ���]-x�c��l�!#��}��� 2�>�E�2�a��=� T��d8��h�����
��F�����qt����%�sY	yY���`C0	����/ �0]z���,�r-g"+=b]�}��孛3,߄yG��x�Pe5�5h[�5�u?�i��敾ȫ�\H�6+��h)x�ߥ����|���`��b��I+t��5̣#�w��V�mi��5�o�Ia����;f=����H�N�4����nܣ-��	USg��9���ć�vژ!#x�d�}o&��h�G/��i�Icf>�տ���O��E���	L�lϑS��1;VN�����-�t��E%)V���Rq�#�wwYZ{�%�x���A ��v�\���#^/<�];��-yZ1��+���/����{LN��=ER&�/�wS��xt:��I���C��TW���`vU��������Iрr�J#�e�ד]��1���
�4}(���R1t7:l��*uMgJ���bX��GoGO��Ņ���06̐��n܍K��nuM���G����҆�J��jq�i7�x����Y�вY�3�c�y�\�f�s@IK�� D����*��u�_A4uӠ��P�#у��f�̶��_����r#��1-L7�?��^DE����3�'�Bڪ��.L��&.�U�C�I2g�d&(I�1�V;��+`��v����38�/=��ƅ��c)�\ϓ�w�-�`��]p�u�n�m�FI��B+�7jc��P�>�b�B�1E����U��J�,}��Z��eb�6���h�[�-l�	���s,��E�hs��E��ïkk��;|��F�;X"?L�hO��.����?g
�Ϲ�! ��j���\�kFR	�c/��z�j��8�>w�9iܡ�����.�_�� kg�T���;k?�ՠ�ቌĸ(۝,�#Ve���p���D�v�$*m9�.p 
$�$�,PŽNo��P����
An��7t_�n�GO�Ѷ��"��|�^��z�蒮0I���Fi��\�m �M�J��;�/����F1{�~�Uk$���#C��y�;^:f��"��`ۣ�������m��&\��p��G�_/�ҩ�3�Q��9t�Î��dy�s������0���&�y�:��Le��U;=è�Qn_�. -���Әc���a����r��l���\��;ެ$] �>I����w�:C@��Iers55��0]�&4�d�Aݜ����L����
�[¥s��5�V����H��0P��>>�� =?���m ��\�v n#1��j��S�HLN���M�R�^�[��4}@.M�	4U���y =��M���M.���&�TW�8vUE�F��ʖY�$�VV���N�'��@�;mQ������˛�?ET':�&Iz=�U�.�󦆯�!��K�dG`�>ƾ�7W�;"����i��<	z��.��V�y��]�>+�@o�$R"�p5K�� /��h����,��+�ѷ��P��m�$���C�����\�0�y�]��u��w�#�[�^��F��#Uq%�}���4n�3�*�N�����V�����~�� )Q�yA����Ɲ1��Yx�����wO�� n��T�[yY_b��tt����M��R������A�����ul�Ȧ��Y�[OD�:z��4D��=�{3Xg��e�ş������ҏp��]�ɴ��"�ܪ��e�˯���P.Y��[�C�_�t)�Y�����b��q�߉�����	<�������3�S:0M����9? X�)F���j�� ����)����b���GNb�Kߎ�%1���L��X�ѽ B�T���Qm�u�%��k���YV˒���;=�Qwѱ�<��$�n�������A���Ύ�����6���b�Zd��^l/?��f�P��e`�9E�����4�E���xu���(��ؙ��5~C��[0D-%_��o��w�h�$�cj������b�ڠ�Pn�Q1!ɕW�,��$-�Ww	S�r��X�}
�{\����T�D�t�B_e
/!o���$m��4�ln���2Z��k
6���Tļ�Įۺ�>��B耓���-������@����(7�:^q��K�XH����ul�j�R�r ˴�sZ0���(�:cg����@@ٯꟹ��1���l��7�F�����r�u�H�s�um#��29�����*v#��e ל'9�N	f\d4[��{`��U���� ��Z�9,��\�R+��2�H61�t��y���(�1�P�d���n�NY���p�oF�Y����#��G�Dd��j~]U��Kd��&�ϬA,��]��5�E�G:�F�_-Uڗz����{�L���㛇��(��-SOLCέ��km�өG�B�V�F�3w��N-���([�1�h���YZI��0\���������r^q^j���	����"�x(�^�(��BQ��:\~6ߨr�5.�����6;<�q6J¤��>�E�e���Na����߶���;�"�N�v����M��Ժ=D�8�E>���4YJM���{瘘iP[���p� ����`��U�� }�"ۡm���%��c�_��״O����^]�\D<N�#m�sPS7�eRvt�7���Tcj⨮��<��î��xe��(��Ӫ��Vz>JC��m�>�kl��0r����
�.��@s5�bL|�`Ԫ�i&�ӯ��}��cpteD:��.��q+Ԡ>W엃Z���"�\���!Aݤ���u�%�$9�põ���3dH��E���(�A���6k�m���_)l-��D(��������Ӯ��.��t��/`�rL;QL�q�S�kTRO}[�N�W4�8&0���R�vv����<3�������$�p���CPLC���p�������3��Q��]����tV̹Q�E���6p���������Vi^����+i;5�Y'�LL➂=Y���ذv=c��������Xxd�����J[��9Te+#$CÀ���G�Ҭ�(��V��d�:��,'��׳Jօ #���,� ��ٮh%�Xm���?�NR=��g_���7�[ $� ��80L��/�(M��O�9L��i2�QL#R8Q]ܻk�}$��/�F���$��
��K�BS2��0ۺ���w�����a	�A�o���$��"|J�W�L���g��]��$�WH��6�#e��G/7ؗ�P��㠹�N3��)�&��
C�8�\�(:�y<� ��Z��	3L��A�������s�>��;P�����~��8�W�҂R��/8� Nu������V�5;���b��m��6΄�:���</���`���Z�*S��zɥ��a�@�a�T|a0Wa��n@���oY�G$n��1����"�'�XX�_���;��SØ�g+���!#�Y�[Aڶ7�Nrcj�D�����2p��q�S e<��^q� ,T��.����1�n5�>��g}'r�n��2Tf����-���`���YS�&�붛Y8�7P�^�ds�PV���g>�+@�\� /cc�a�����#ZN0�;���t�]�7��O-҂8��]l/GM+�m+��n�안��l��Q��z-D ����m�T��:���~���Pg0rL�V����B���}�Vu�X{����y���D����C�6Gv��,j�ڒ�V��
����(`~���b���bfs�[IVR��I��&����vb�,���� �п2	}]y�AY��ApM��(�;�;�4����c=r�z�n��
���)E_Ä��F���g͢1{Y��u!>�~��KZ��������,z�f?h\�__�6Sj/��&?�Bٜ��u�dNb�r�9d�����k���aAc��D6CA������y%J������������? H��L��������y�hj
��M�L�O�X��vd�/�b*���P#n����q���|�5*����w���~n�R�i�j��Yh��x�J�G�Sm�b�]u&�������N�l��f����|G��C�u]xlծb�Z��1%Gd���вꤐ�ۡ�Lͺ*a�R`����)�$�|���
B���!5#�Eo�+!�*��)=�m��8}�df*��Ŀȅ��EO�x�4;۰;�[�����3�1)��E �h�G�g��(��{�k�V�o (�n|�i���MfP��e,0{�Zw���C���A�b��1-ދ��֮����[�[9N�Ќ�9�/؊kK(�,��ͪ��Az@���o��ר3G��ެeT�'Z�����C�(Hy&�aqqh�0��k��!�̠�ZR;.M@0I��r<)��τa&}	�^�a DE)2M�2��Wi`.��:Y�4�IrWb��������:D���>������6�����*�4���iW�v
>ye�=�q,)��%���U^c+\dY��^ꮈ�ߡɫ�4r����k�dD:%�BR>��G��y����Gq�������7q6����b��R*-&� B�&���� İa�y5�ܝ�5�uΝ]Mưހ�ڔ��ڤ�1�_&��Ȓ<EDml�Tڅ�h䘓�q%[��;�v���x��3au 9�IK	�Q��_=�u�,�J!U'�ڔe�.-yR*t��A^,���Â{EܞRڐ�?up��>;k/��D���B�\\� ��~�0R0�� �E�w�@P�ki�RXs�гx/ҾL!������]� "����� Y�;���*�[�&�������L����M��N�I�H��q ��6��y�x!��u��3{F��$��]�j��Ӫ���� y���f]b��ҦZ�u���k����8bc�M���g��Q��}R�W�{�^Y�)��pM0�B�F�+XA{U�8t����eM�W������_(��Ls��e0	#"IbKjǩH�3�1&�c�0*�e�kF%����]�gB9����Q����j���3��EٗV͜�g��z��;r��
303%�����}4w�M���d�!� �&bWh{�+8e�G��A�,h��^I	�]�����^�e3d��g�	4����c���y� "�����=����	{d�����/q���O��w)9�6�7��7&���;3�H)��J«��tR���O5?i���ȩ;��7��d�+�Q�����Z��z���ơ��⛔Y�4�
Y�E�4	�\�V�%�q�O��"���t���P�/S�eإ��х܏u$d2���z��f"نD�3��p��rݚL���;�v�ψ~�yo~k���n����cQ���+��O}P�I\�P0�1�|n��vI<l�����D�Z�ڇ�%�ڿ	��QS��p�8+6�2O�"TW��u;�Rh]VK/��,��ڢq���p���p�c��k�ٶ$�u-(��c^B�o�2��x����3�CIWvY���
F&����X��f�[��w�I|QI7�e�g��s鎔�]k��ε��aʮ��=�(%���9��
��Uӧ�P'�r}e�̿T�LUr�E��	1<J�'_�#���6d+�`��.M�/�w��æ+�Bw�,UT�5�$��L�w:�t���:F5�q���=�U��Bs��胲�f����y��ܬ4+*;/��P�9��d���zu��.xQ��yZ_��zt���
+�@B���Y�x?���p�6�^��YtL��T���jJg<�KT�k~�_���5��i��P�v<�	�sSk:��������l���㥮Ģ�q�+��1�.�2����2BO�}�t�6h�`�T'0���!��}8��$�0bt"�jWb�ˏ���v�a�pT�V3Us��9��f>�7�Q��E�1j���{��RԹX6��,"�򧜖L���nm4/VP�Ob�w�CSy�����k6daO�1'ue��
��چ,�:�7o�:9'/_���K0�����%�PtNړV{B�M�]zX��N3* z��C�&. 雺��CK��Y��g�?���U�J��W;&�z��8|qj�7��c�h��B�m[���BB�Kۖ|-݀�Ģ�>�s�g�b��6@�*�Ԥ�ɖ#7����̷�Ik��Ve�i�s
sG+�����+u�� m�F��J�M6y����Y��[a�
��
L���{Re�y]~��-���]u4M�Ю���:2�U�����)y4�v�<cj����`X�4�Y��V׼K�`9��a�e����=�0$��@� ��I��m= ��g4r&f�N[)��?�w/�)sY��C.�\Ʈy:Ӿd�$!�n���)	Q�����u(*R04��:���؄̈́͢J��CZwm��g�
����s5�a�i�`K�N��N<zJT��񺫈,��lxO�#&���`��Wj�k�l@��E�b�6Q���G
Z��rP�h�O��D���L��-3��	R��v��� ���d����#nD� ����Ie@(u���r"M'&^���X��$��]��3�z7a���_Gj"�Y�t~Ǽ�|�	���qp��C�Fj��QPgSӋ�p�O^��]�C�������t҆�q��A��\����ö���fA����i���$����  	c�%i��a�o�q�Z��_�Bv�F�..2L��R�w��� �(�����jr�W�=;�����_�{�BK��-%�ש;�%r��+`�������k_���T&P���=c怞�*�_v�/�V�~�)y_��u�o�A���$��+i�z��R��I�=@S^�v��b
X��X�肦?TٶZB��ɭ���j���vZ�{�C_r(�Ϥ(LmQٖ���E9!��,O+�<�HxeX瀇�����V��O����j�k` ���az�*��gωc�t�(?�<��
�G;�#ݲ����|[��3�NxWt���"<nW}��+.�ԍ�x/.�5� �&z�&��E�E�(������A��y|�n��~�*Q�s}4t��>���p�1AK:{������EE~�R�������}:��(Ay^6'��� %����l^l�ϡ����o�~g�F�ݗNS��Rb�潤�{p9:X?
$1�Î����B>����X�Yy�SV�QI!�s@���f����!OQjмH����]�k��#3/�y�cb�}�oxM 	ch���NvDَ���C^Lo-sl�g�"f�����(���� ޴m��W�P)��kc�m�q�g쭦g'�ڭ�`z�����)������9U|e5f3�|��&S�m �4Y{,7��J-���p\G�	�p�����A��`��:J� �4ttG\nv��h���K��C�ʯ2xm��-��N���i2���՛�#��Á����m5L*���aW�N��{Ύ���D�8m]K���nf�n+�hv�^�/K�FB�_��� ��g��U�u#j�ϜT��U�úӎ:������P��d���jn�:&��[��Zѷ�Y��j:#b-�����Ni��_m�-H�ޔ`�t���ǋ�^Md�ϡ�]�^Sپ����W�.�J��(�/ǠǚI\E3���{���
f�)��0�k�~�\,� �h"�b�f>��������ճ��g���1D�5��Y�͕�
�]dG:�(��%3	��\j��fKp��x5�/�ϧ�o�I�L�ųYM�L����(�Q�|Fa�b �9�:�(L;K:�b�%,��d����n���]}�1c��FO�(؏�D�����v��Y��Ӆ�H���@��H��w ��tC���O�ȴt�0�����}�B��`<G�EUHi��8_R�0���pd�^�����u�;*J)�b-�&��
 I�g|	���˂�����:=&N_f*U��m��O�%����x�S����oT�+M��؆Tx�C��;�d�/���26*#f���P
NF4��{��U��a��k	ʌ��,���+L��[��q��I�P����(q���Jɛ�Ά��5eJ�^Z�*f����-h(7�y�9���L�?��^8� Czd�s�q��P4	$3�+�7O��o����|� �H ����k4+^쫇���Wezi	�<i��2>t�M���w�Z;!��L�~ɆS">q��8����x���U�,.��hS9 ݋9�lH:຅�Rx	$��b�AD��nɂ<z�P�����	`BJ��5��pk�I+)��৶�.�[��e�w:>���q��r�;vH`�Y)]�S�b5SB�� *���{b%ŦU�G��̢�`�4�9ve���{�O�g#֟��J@�R��Q7�H}�U�Vz�!l�v$���]�\���-�)�sq��X̮��v�8
.��,`��[jC�C�X�ת
�C{lZ�5>
6	y�6L(��;����D'������
�x�_�m�{j��W��+�i��R)�>�)�b�d���N��;�v_��x�g(�!? �RW��t���^%�1 ��2�L�r�����KθǇ�=r����ҰzȬ����T~�G^��i�JM�����]D�/�t�듯E��X�musZ�*���11&����D�}-5I�ﭑ���e�a�6~�~�U�܀�kwoxksrq�'p�Wm�qXH�i�Ƴ��b����G�P	܌\��ۚ�4t�ٺ)��"���F��RL��5�<�2�9o����&�^�(4�q?LH�TE�@��_���	��ܦ�)�7�a ���k� D+uI�or�  8�6&��^��W���ɠ�C��R5iҜT/��3�y����>�yy�aYoւ|(�19�k)���V�x:���x��0��#��og���޸��"vhC�O,R�}�I�(.�tn�pٸ�t}<��e2/ G:R�t2��;��� Lz	��H�u!�9�y�m"�MЃN�����؀( f�a/�.FB���P���nK*�މ�@���C�Z�w�V:9CFYS�R��L�pev��z!i��l̕ ���#��jҧ�hu�6��n�)�mFA���3�_b�4E(�&�����3�fs�͜��P�z.j���"Y�yh�T��q$V2�֚�I�u?�����e��#L
8
A�{r�d&�>\��wV��;ۇ�=Dz��ݹ����&��#����� 4��f�>Z!qr�����49a&�]��/0��)�������5�7�5��5lB�ՆS��v�_hՠ�K��q[�	�Q���l�`�� �Y&���l����hY6ܡ{��]�6A����'�/I�/@j����-�p_/K�ǯ�/��Zbp #>���X+��A>b����m��A�P��^�i�L�BW��xr�n%/+��E ���5"�,�f��C��'���Ph�%�6��� �����mii�����5��{��,�j�M�|Z��n���������fe�[���J��H�u@�2�?��a�K-���2���ʏ�nd�A�����J���}��ȕܞbÆ�dX�!���`���c���/�x��_L�Q=+;;�)�7��zu���� _��5�@2!���Ǩ@#�Ô�
��a�w�\�"��I��Vb�c�-/�-�	֏j��[��/
�o��l��`�p��b�]��?��"�U����9�^��Vy�L�6I� "?�<�`S	�cZ�Y27q���.T�e�ѿO�xG���.�Y	"�鬵���b���L��{.���M��}$��!+X]��eiO�͌����U���H�G���M��
pĎ��7�NT�,�ܭ�KD�����#X��;������u�X�@���#@�[�Ku��숭'!λ����{e~�B���-^�)��ʜrN�����49��6&��#m���{�gi�m�Q�#c�S��n{�H"�B^,�ˌ�z�Z��(���M<2���3��õһ�MT>�S��8��F����8���'�Z|7�:�Xw�\�w0�co?�*�ij����"q������'�����p��^t�??�u\vĴ:܀e���2��z�L�<�3����l��褡�!L���V�^�zѐ��7pd�1����+�]��>����A�t��`���.��H�7��B'��/KfG2�뛷7>�;��vk%[�2ȝS��lϤ��E0c*��R������Ē��ȯl��XSrk2u�m�謑C���AY�Μ
e,#H�B��u&���y�A.��=��IK��p��썏�XQ�U� -�$��g_�}���T�t�
1��a����>?~������g!#^��I���P	L�|?Gv|N�5��A� ��/��$�n�v��o����K��i���1��Ĥ����#d����?V���M��U�d((�5�n�GaD�>���c�pjR�X4}�:�����m-�O`y�QA�_�o�VP��~��6e#�HҌ)��fZ}���
�+�����9CU�~��Q'�n�,Ym��2��ڄ��	J���2~(����J�S����H��#�$�j��9�W#6�Z��9I.���ۮ3Ҡ����&�"1�͒��`�>y�]���S+b>E�9�z.�h�iBRʪ��ӬiԗEϚ���1Z�k��F��*�y��p,䞄�������-�!��r�70^�cK�-�h{Jp�Ճ���$�εM�z�@��u�f���h:�L�C����	Ǝ��Nt�A}a����������Mۖ��QӚw�`�%�[d��_5�fҲ36~�	H&����tѶ��/՟e��MIP�S���n�$�-3e�;N��P��I���ݰ��KE����ymJ2�����>�����b�x��j�H�B�"L�*<sM>�y Η�L���NH�P2�e�7�ciqi�ayg	�Q��m� зA5`�w:�O�RǪ�s�j\{���ދ_�;ۼ���W��q���U����W���J;�z'��q�I{�j<[엱�Ï���mc�� V�[�S�\'9<�>�����ЎK�A�q�7�b��нuzb�v�q��U��!����C4��tsd{ߋM�y����@2���sBi�4i�{:��e�b�Mũ�-ɫE���iꊏAT�;p�y����9vo̭mz���3��]Y!�D�'��������Z�	5p7!�G����Mį��-߀&2������e����LړBWc�s�&�_n�[��Q�W�Վc���z�~x���!hu��]h��ⷡ��Wl��YB���LƳOj��[e:ze_'������4)K^�AO��F�D�;����޹�j\��cￒ �\+3����ytp�c��0�Dl]���#oBX���D �N�Y��Ӊ�~ʽ���AO�?S���E/ae!fgYe�����H4�'Z["��V�t2��x����\��lP�H�����w'> ��J����3,�e(�!i�+Er�0���UW�˃��P��i& 0���y�a��W��a���#V~׆� \���O��a!�����x��ǿ�������_@��)���:ɞ
u����Σ�ʲ최�ץ"�e���^i��W�E�9��'j���lk���++G��+����4��E���t��m���3�b"������#t PWͬ����@�!h]� ��0���[����'����ƿ�9#D�H��1k�����Oƕ%�Ȫ`��*�ny�M��Ө���4�V��h"BL"�1#��4ù���Dd"_|���N`S��'k��q��ݟ������J6ϯ|�Rڂ�E�}�c� 1HEgv5 #2���r����ӑ_�}��Ӯ�'���,��Y�Ӟ$�ۿc��_�;_��@r�ז̼��u���J��L�>G��r�M9dz�'���N'��&=�&�#�jƍ�5����x���щk{���Rp�W ���Ͻ/E��v��A�%�I(�n�Mz�w�X��ARk�/-���z`�c��l(ך�����7�FYT��ϧ; R�Z,�<�������-��ec�Y�Bm�l�<�A�1�v�J�҇�t����a���w6�E��n���@5�߻U}^���*�� z3�v,�v�1���P���� s�h^(s�w�M/���+7���'Q`1�)K.D�L���.q�,tlD������n��=K���k�D@�~\��������03SM��gTh=E��gk�b����M�����$I$���㣘��vHg{��}\0��q�z�gۏ� V�#@^��Eby�	��u�[����l[��t�M]��D��������iKEj�|&���ǐ�S�~Ҽ-�'�ʪ�،�����-�V2�W����ߧTx�v�����۩��{՘���K��8b8�����"�?�$��P�a7�6�ч�NE�0���^�j´��!��2~�Ais��_r��F�ڜ��-b�$�Cr+�벂�涞l�6��2C;� #:��a�4�|��@������n쉪����c�T�҅�e)����Q��$dh�3|��`�<I�Ĝ	�x�ИaJ�3�á�^��Hpߥ�[��' f�S����u�xB�jP���s O���m�Ȝ4+�+���b�Tp�m��)��`��\`��5)^Z��(.I�4�&e�^��HAnK����J���ǃ��/r
�8�fiux�X��}U��}[⳼Bu¤�\����"F���z3/�^?���W̿�#gd��{h���˒�*G�9S6n^�;�jl������ܬ�-��)�YD����5��9_��A0��AR%n,��:��t�A�6nM�-��:^��o��j�.�>2MjPǗ*�:�^u�l:����s;��]�U��e��P!a���$u�V���FH�B�y�TKN�� S��nV���&�A����8MK��e���J�`t������..�jA��5��o������-�eM����N�C%Zа�I�3ek����Ο,�'�^�%�)*H�3lJ�W"�w���~g��(--��$>e%gF�����ʗ�h��}-��7��N�$����h̢��rB�{Ta�ljp�!P@Y�lIS"�x7���B �Ӂ�e��IO�����}��PP+���ݠ�V���9\f�ƎC{v|m
Խ�m`�i"����I�rf�
VA�m��d�7�����w�" ,��띍1�9��9�-��ѳ�0�j�F��=`�$|<�w�����e���
��o֠T�TO햸���� l�0)�[UےuRN?�!~��e��\<����a�NQ���[M��>iж\u��������p)� ����GH�+�ՠ	�稸�TGͿoh�I�V�L�2(��)��,�����m�+��I6A�4�˂]u�ix��w��i]�e2&�B��c �<�5�����n�&�d�NwJ����NUQ3nV�(Dĕ���8�^�余@�4�>:��	f�:7�i�!�ߣ��؆��P���nv!�>J�.�����!nP�Ą��V�@����6@�1���mUa���� V�IO�,5 ���k��\���?D�I<Ie���-��]�]G��,G�6���氜��:�o�s3'%�����8��-R�\����31��q����a}<O.>h�b�v���Q����ȃ=�'�����o0Â~�'5��{0T�HOOIZ�2�D���6 |cz��.����L;~4u���痃���k�N~�1�I�&@OƗ8I�8g���]���2 ��#
_Ɲ���M����r�?�_7s)��L�h?<Hi�������Ν��b�w��$��ڡ�ۅ)L�^x3b&�&?��}~1խ�?�S�J;!"]��P�_R�@�B,�A�S�u�h��-�X>W�VD/�q���+���C�؛���~��cz	��7n�ݿ�!N�+':�3��W���N�J�?`����Vt��~�y�M9=��_l���Eه�Hd�=ޒ�� �|���2c�{��{�*�q7;�Ie�2x��!<ojs&Q\�?ؓ��n]z\��r�p��C��c`����Uc�7i�8 �d���ۊ@T�E��4+�c6��5� 8n���|�&ɷ��>^��t�*�?�k���w�E�X];���Et��u�^\j�)?�ɦ;~��Ġs�JQ#�n�JBZ�u�C"O��t�P}��TaB�2y|�q��p��+�eo���Tn%·ө�??��(q�bҧɉ�!�_)��K���<}���h� �P�����&��MϋF8�	+����	�<��R�P�'D+�d�>!�p�
�㛴@`n���{�+k�C&"yj��;w�Ҽ�5H������~P4�E��ᏦO���x n~E�������	ӍZk��F�m���¯"���W+yl#�ep�`$N̊���r�u���b����-zN�$a�A%{(�݈������j/��z��wIf�QԫЮ��񓫽�fEш�3z`��sf�JFszǑ�ܹ9��8��%���&�,����<��E��G�N�����sł��Mb�ʯ�l���?�(I�v���}���^#7�}J\�p�>��^Of�5R����/����l#��)�9[G���0� TZMH��xe�]~��B��<�qx)Z��t�E�ɽ)�)���0R� ~����(�2b$q�΢!�`�=�}ѽ^��U�z;Q���ߴI���,���/N8i��Y��e.b�n��*�#h�=HPR�{�����|Xo(e�:��;O�K;p�V���X���u�e�d���Y^���#ѽ���ӕ�o��iD/�;wv%��O��ji�m�dPv������ ƀN�>Ic�-�;��E����ǳ�t�s�/�zJ.Ŏ.�VC.�I��QkG)�B7�O�X��a��e���(2M��}�cωc�>y۪�cUn�[i~x�yCe�ku��箼����D�m�VT��]�p�ή��F;e��0�	U�1⻰A�H@D�o(*۽y]��t��&�"����%��hqS؍�=���sY~�sV�1��m��5������O\x�%��6��P\��ߧ�V���X�m��k�^��ߘ�Z��t�%�lݖ
K������
���t���c�*����L�z�`Ԣ��~V�K9x�-����5������e�i�ۀ�ٷ�V��C~���0���v�F���]H&!�*"Da�6|'����zѾE9ģr��^�Ֆ(�༶$������a�l�1A��a���Ʌ�s���%_�
�fS-��lC*3F'� �j���
j����{�OΗ��?��� �s�P�Ț�ӭmS���$�a�4I8���'�J{cF/�z�4����h�*$ږ+xl!6�����J��[�7�N�5��{��%��1��`Vf:�)�x�<[t�8��g)�~\�5C���
��j���f��*ʅ��dt�#�"淛��4z�VN�F���`�(�V�a�[���$��̙,'��#N�C����X�{�P���>���V���F�YA,Z���������a-�-��Lլ#�(�b�O�x+0]��۬(1����?�&�W�]�Zc��eYʵBak�ӛ�8�zR���⥢�J�pD���xU%��Go��NrG�r�/SX�w���7�f�]U᥌Z3.��9��r
��
�8�Qq}�I�f�0��/�w��?L }f�o7%	�U!��� WUtU���]�[�,M�`���/�;���_�>6_��%3�cΣ]�0k�W+䂔�.
�W��fY�w]��W�A�SH�.�>�Q�"Øᵩ;��f7���9�ď�N��JW����3锝���cl3���5�}�J{�U���K�B�a�5,��6�؄�S�L�pO�wvk�hM���y(��R�у�-M<��7P����ߴ������.�5�����)�i��R�׭����7�
Iۑ����&{��3`�D�s���U��ϵ�O���|����SdPW��B
6�dz����������\*`Hc@Ʌ���"3P/ �&��q��&�����xu#'�}�=$�b�v��f�\�3k!�\o!I\�N�^�p"2�vU�=��&��{��<��8±��kw���?��eE�0�c@ ��,Ӭ��)���>�w:S7�����ˌ�&U�|���u����c�Z�':�;��}��&-���麏Gh��(5B�S��V(Q(�:e�b���Xx�?�%D?cVQ���&�z8M����RE�Z"F$y�%�h�*>+��r�p6=���1y�w�C� �REktKp!��=Aڹ�fD�Sp�-!*0tFyF1�5�QW��M��2��?������`̷�a�����( ��4}�Dpe.���4K��o���[��(NO#�tx����#7`*"�m(�xl_�?����d���dC&��qNB/��Jqc�'����>�Z�C�g�Y�|�~J_Qr�@=�:�a�7�Y�%o�Iu]K5��ׯ%Nk-Ag�u>��t`M��{Q�-�)�{�_Ԩ�9Y�ǜ|G�$�D_�~����/��XEw}�}X_�yͽ�5� �e���$\	�S� B#�~�cH��v5���O�4��a������w��MCtج���M@f|r�������U�g�8	�Sn��&��,�v��g7�,�*�@��k�^�z$�DvR�d���K�C�&	�,��8�uJ�y��Y�/�"��!���CO<�����g���cQ.���5D\��������z��� �#N�s Z��Y{���"Phs>Yw��Y�t麦��Ʈ�ِJ.����,Z"c
X�u'g�"hAQ��_z��;+�rT!�����c�5�b}^�5T-�d8���ˋ|��I2B3}d�w�6���3b[%�����4��ߜ�UP9J)��N����3d�%}����eO0=Vg�E_������/��a�5�(�)��ƺ��ߔ�a����-��}�r�bs�U�݁0�y,����/��.��g�²�5O�$f�Kb�^'��]�N��GH.�t!��5DIE�`ס�SA�������W@Z'��Y�@sX�}S�R���:�+4�n��:%��Y*鴍��H!��U�Y�X(�t�`�L�8
i�\W��;�JV��R�:�k����:̼��ɈLw�	��ߘ4�6�)�b���Yd	��|�N�?t�ge}�lQ�T�J���t,*�[�ti����8��!6�|=�``�r؉n�AHǻ��B⭍2L.<9u!A��b���hru�7ײ9�c���w��E9�;�" ��o�3�d�7~�F��� 3�gqhHG�M��$9���!��/�ƒ�S��%Q�#���N.�Ђ��2����ЖU-׍r7��D��>�ᄒE�*B�F�,٪��4����h'�gUf�%�᪥�	�9ݐB7c/�-N Td߫��\4������>	j��A� j%�z{��%��?���Č��Sk����B8�z��w�6D�D0�`"_^�m��"�h���F����9f]�5�����A�q
;�� 0�`��E�k��_KR�M
v�)ܴ�i����鰎M�c�'�R��~ڞ))�:��C�"����ק������X��E`�������]�q��(A@a�V��4c%~�8b�`B��#pj���׿�*6��	6S�L94�Ļ�ױ��y �]A���{���	8�Ba�����4�X�u�!��z�V���(���f������ׅ�BƜA؄�4���y�	�e��[Vk��&ry��'�����]�-�%�J�$ h;r���R�Ƣ�@��S��-C�����0)_���]3�mM�aM�{Y�R2?VB�����SC^��$b���?���^�����3�)���S闐ӑ���-t�$��Ï&8am;��*��58b����	��o��b�Σ���#�����44�VV� �ZҜ����^�ζК<c�u��1	2��(ꐢ��P�mB..+�w�`K�c�^�$%��,�ٷ����0q>S�1��t�+gI,$��18�m����d�"��e'^��d���e�}P{8e)�~��Vп���Ձ�L#1��e�e,?f�G'R�F��u����/�m�D�48JUB� :�����;����Ek���q�B��oG�KȈK'�Q��Q�/��sRd�Ati��%XsH@b���<:L�ӷ�s�s6��B#czֻH��cFP��]��58�ȕ�p�YK�f[��C<J���h^1�����b��г��aF{G��E��S�
yW��l~N��qۂA~�o�����o􅥝�$R�l�F�&�qƴG�o�#΃�>v��z�ܾ�x�LY�k��?�ra#�"���-��Mu}I�R�!�MV�"�+�T��`���s`c�1�I7��xQ��.\�E�Bd5�l)u���"O�����SG,�Y`���V	%���k����Q�����S���daZ��
�I�S��&��m�Z[�ƾLj"9xs��{x,h��7��9#���J��S��	�K??��G9^��	�
ӫi�L�Lb�.�5a�aޯz��~��Z��yQC��<X�c����I	;������Y�F�\�C�m�[�i�d%`aL�<� 5����Tq�cp9ctM�/v��I��>m�(\ i^�)X?<Pd���G�>Q����#���-D��SC:�ɚ�0;���!*SIu��o�������5���̲���NA��;��Ό� ��SaLH���1>7�Lr�!)�k����+��	jИ+�5,Љ�Y	��m� ���ظ�2�ߗ����%��yۢ~%���b��:� |Tϑ�������d�$��O��K��j�-c�"��P��������z
hn�7Ņk>�+I��VS��e�1�-���M��TįŤ�� 9�쇆E��{��؞��.�dB]�27�y���}I#��?�um�Y5Z~��g��`̥Զx���I���1��Lr2{ƹ�=���"��W��}Y<�����	�]��j�NB�jzq�c]����\w\*��<�������)$�<M�f(ш�h�|:'fC��ka�}RS�2���A���B ~�����ce��I~�ƛn�9�۹	&��(��pkp�z���&�C(��+2���B�l�U�����:�6����VM~濐��h�7�$����S������%�K��:� ��"5���g����ԡ�g"�bSQ�2�B�� ��z�P�wh��O1LC�es�`�k�������l/T0�7X�$��b£��!p����ϥ�~ۗ��Qd7� �sO��6A�՘x�H�r�3م��v8*.�^8%G��u���0t4��z���q� �?�i"��T��{�q�AΕh5�'��O�?�B���ou�A�'�5 k�Z��������B�D�N<e:�*��*�"�!�)䬟1T���6��#;L�]�$��5��yz'�ŹF�7�u�W���a=��Z��/�̦��&X���Cn.c�� �Ϸ��ړl����O:�`�g���k"�W�����E���r��U�nv��`���|`��U�ٮq>�[�~�4*V	�χ���N�=Yj*c�~��{Y������r�Y_.\fY�{��U�H�$Q30��x%��=N�FDǵ"M�2��:	w�&��bD��x� �E�_�� ���Av�Š�4���=��m�}�.>X�RƂ1��^ŷ�sC�Z��@�(f�^tlߗ@�)��V�*���ۛN�:l�-m\_����iuO*��m�p�����\�4�g�eO$��Z���>�Ex�
�7Z �����R�|� ���TK�t�(��WMܧ�[L��?��qz{��*&$@�e)�.D����.w�|@�k#��q�`�%�~`����� \�]=��؝���ʰ|�ٱݺz���П❯��SI�}ڀ��G������2�(гp�%�7�l1aޣc_�y�yY���>,��8������� �v�-��D�w�:T��r��r�O��['��lӊ600��exLf݆O�bRB��gL��zi�c%)�ÆfTB�#��Y�㎾Tl��^\�L0���Y�Eu%�&@����\zjZ�:7�����X��y��|M�S6EC��B�s�\-/t��\Z9wɚzW�>�(�d��:Z�����L���ԣq��)�=�s
f���������T�`Ar��ץ�A��8~L���uS�#E�Y�i��+�@)z��?<Ց�G+�^�D!L�K�>�0�H����8%e{"����3�<phbq�,�Z���A�%��"и�44���u��10��� �d�\=�M�Jur���g���xH��4q�����ן��w4h�|c
��MV��D�F��B��t��oKd����V��͈��b����o2���0(8Z�z�?���<�� ~j��7��\}��]�ح��w�C9�,��E=(��FO� �.�5���*����s����_]۲�ϴj���76��bb�</���`$Л�����j�W]�^w��+.�� �!�F�m���|��Wɝ���˙��W����w�q�_R��
D�UJ>��ݾ�|�:�a�Q�3^�=8󿀚���Fm��)D���P��8`r�F����f&fO��6�t,UXd��/���k�vO;e�W�?���JvR��E�C�{9����~�BT�▿��G;/C!`X����?�6���_��s۰�'4S�ч��_�c���Z��GMy,@,�˿���0��Y�8I�:R���Z���Ky3�G�n�������$��@Ǫ�����(��	\�����/LA&ە N��kK��8l/�=߂�܈��y�f�IT���ġWu�_Ѳ��};A��~�tDs��4E�{��G����Xh�L����}�u'Hl {�^��l�I�]�gQ`��_3���e��'��[�T����ۼ���_�/��qe)as{!%gb��go����Q)VFE��#�-��Xʢ �P褘c�l��g�:~�"�[��?K�̽�ټ��eF�Ci��Q�Ĉ�Z�@�8��^o��C��6oy6"��T��mA�#���B��"7Mr9 ��$���}� L����BTa�'��6y�L61���+385I>6�O˾}��x��f�1��f%-Y�@�j����;�c���z�E�?R(5_�hL�da����k�_/���b;��֌%+�@����itX��M�o�3��~�������p8$�W �ɸf	ҏI��-n��]+(��:�Բ�~Zc75L ��n�1�j��5�吖>�7�M��XJ֢^���(wg貢D���-CP��Y`�u�(�H���J�cRo%Ӷx�a���@}��m^%ۼ+1|r���L��!"�Tӧ��X"��yg~��5Sr���[�JPXy*��i�?PUz�r��դ@5��4U��t����Kڽ�_��{ /��us觠ɯ~��� �Rkͯ��K`�e��hp�����hk�و���m�I�/���I��q^�������U�*g|7��0ST���LR��u\z�Z�# "��|d���sYXrBe�ǹ¬�����u�dӫQFm�M����%~[�C���N���c������)���K_�JTλ��u�g޷>/��^{>c��I0A5�뱱;5���.?�I�Jd��hcׅ�u/I�'�*��ӟ�t��̎~��W���T���llR��)I#�'��d�3{�oNݗα��br��$������k�ɤ6�!�>�����x֯�7��DQ�:T2�$\헡�& T�K�^l���rqh��6�A�.kTļ�>=5'1V��o����9��x`8�}d��>~��f�aG�o鈤=lф[d^���sn �H�u��Ǡt+��ƏE�]��"��<�����4S�Qh09;"�H�kM+�0�f�g��n1���Q�
��������<�����S�d"�:�\�� z\~ L�h	���u��6I��: ,�l9DU��ŜW��@�L^d�V���l��a�Uf>u`�NbW�A�,�DAg�X-�)[�
X����y�Tp�8�B������4g����IYV�Z�����%��k�H��-�]��jXS�'x �S��W�A�FA���Y�S��}J�ˇ�^���&���x��lP= ;moe�!���Ũ����e����PՠA���`)Q�u���J��M��kEtۡ8�����Բ�Àl1�Y���fˠ(��y��q�v�P[�v�����x"�.aIG�L3�����{����l���\�~^mln�3Dsל4�! ��@d�uURC��g�S��cQh��<�덄Hא���<|�T�L��"%V�UP �H�̕��Ĺ��a�7~�0�B*�(��k~V���ڭ� �\{�l�di��R���Όs4�zh'�h!$*��U�k1{��h���:Y7����SC-
<�B�Ց�w��T	/k����B`&KTk鹒da@�)�~��O�GRW`��s�u�"ʒ��9Ψ�z&q�S�sPq�0X��()�Ce�ud�k�|_�����֨XG����d�/�bP��}ۡäh£��'��J�S}��0dk�d�Z1� �\��o�.��n*>+��,ծ�sV¹J1�˶�
���w�
t��V��H<㗀������i�ʹ���f���}����u��Q4Zk�S ^~�o.��I�7�|{���;\���-K�d6$�շ7o��c9˙{��6bj�͛
�L�;=0(A�4�=��d�E83�<��?tU��ȟ�}���*�w]�*L_Κ��у�	7��s<�����-����#�H�Ã��Q�� <��M��7 ����5��P�"{��wP�����������e�i�\��9k1,�Cuo���R�$���݃u��
12���X���ZZ�B1�Lܞ�ͭ;4�QkX��ԟX�7�YVJ����N
��Q�
?/�u��%%��L�Ozf�����Ydsx���IJt�R�x*{�?׎j��������q�y�9%*�ڵG��))�?b�����5���NN1����H뀻�bv-g�}���>���S�Q杸'�w9㮰���چ�R`;:�z��m&e3�6�8�}-[��J�8�}3��U�m��T�Ai�tD8��|�ә��~��IU����˚Ћ�*��U�N���Xd_�v��z�K|\:,�+������~7�<��Rkz��U`�zuf�K�,ֹT����tJ<U�����mi��F��xٖ����I�i	N�i/"f27�M֑�RTr���O�Ui�i�eT�,�V���#:!%e�5|��M�~��e��=�[� ��Ȉ��8��z�:���ak]73����^jv	�A������}������Z�tn;�p��jU��� Imi�5��u�d��l/_Ӟ7��.�xV_�O�2�)G���A
W���U��T���V0ʽ��x�ɧZY:�Wq;�X�a�2�a��,�<y�i2? �p��3&vY0��wVd^�C�&��Ԕ��"M��N�������p^������1I�@�0Z�m�ތ"�oD�ޒ�C��ԧ\�4r6��Z	�i���T;D��������t��E��\G��dfef,���n^F���[��s?SBF�%U�Z�I3���W��A�Lm��T>e��zl�=|Y���z�Sh���8v���čR
4�R�F&��Ȃ���7��������$"������r6͗�����_��҂����r���@�*Y���Ҝz�-�u�#.�U���M�P&��_��Iiq�v�%�v�}�X���������D
U�-�#'�����˘ o��X"�a"��}��kb�dĂRf*rᙆ���|�����J�E���qs�m��-�0�=�{	f:�b��^Z�ӨO���Odެ`�`ePq�����OG�r�D�TvCJ�������D��	����^F�(�����F���s�G""��o�:�� ���R���K�\��Z-���^z#�����-��f{ےF��Տ"��t�lrx^S�G�,4�~��z�a ڐ�x*�yѓ�� ��o�N��m��p/-ȱ� �� �JR��-VK����/Y���	������a�8�A��t���L�J�c�a�{KX�{dr�7�u��Ӛ�j��XN�!��<l�K��|Yu��7��D�	t_!Բ�H@	#-< + �}���g6F��J�-��r%@;�����#�u�B%F��V8���3�I����9�xRc�{���t:�]e|T���Um-�{p�
_�c�S��A�+�<H��sSqо���g鴰��TKV	��l�o;�O�J|N�f��/^"98n/<��r,p�j�A~��r=�����Y�&]�Ǆ�0�I��H���Do6/�POyO�*'��RRDm�3u��m'�OH[�&f�\D�{�j��%�*X=+D��@C���S�V�/�|F
fmP�k�e��ȣ��i0�P$02��0���Z֚WVD! �#��RV�
)m�I]�e"��OS؋�4�Lt�p	��r9�Y���"�dF�O��&X�wԛ�Q}�[M}Zw�9�j�i� �4B��`�f�ꄮ�7Q��=S��b����ẃY��=�V��TR���!G�DZK=��%�����揕ﬡ ��8&�2�^D�>9�֤n��*{�Ј��ȳ$��"һA�P� $�N��-�o*�N�Ϫ��x���l��'4ZW �O��!ƭZs�e��֮��E���Zq)����
)`"�Ƥކ���#csg��@�C��[��4��������[\��XA�8��@���Vׁ��?.b}
��k����Lf1a�o"�V�3��LW'��	������)t��Ժ��@\C�[3�>���NmsF�� *�%�]0�KoL�	@ɜ]�
��5� Ϧ�c����Z�Ӟ��W]�vIw����H�gY��D�A�{lp�z%�ִ�IZʄ��psI�Yv�6y�8>s�[�'��^����*�su�۵��Z'u �+h��:&�R����?��?W$$�:��^�4|E�c��USxG��)��^�Ti&�16�Y����=~��������FX�Z�~�@��jx�G�+�g�=��r�"��ӊ�s�	ZE�O��Bn��s^�6;�
�]s�~���|gn<o��x�(ԟ�&�T�ݒZ�\a��� ���]���9�4���0 R*�b���u�@�F��r��ƥ�9lt|�����'�� �L�TY�T�[�	�[�D�;'E�����p{�e9Gt�жlI�>M 2l�U�b�6b����L��m��#���&�LQ��;�͐����U#A`�$�b��[�2�e�uWIaA����&r׺��-;��CT��+��^6�(�2ڙ�J;���ya �Z ����$q�T��GٝvQl$��~SТ�3K��Hܬ^m�J&��T8��9����V)/��u�S'	�Sf�1��h���vT<+����F�K������SL������7]�ؚ���G�|74���F���W�W7��\���\d�_58<�Jp*2���1x���L\;��^J���=B8�\)Mqx��3��k�G8�Iq�7O�{�v�ڳ�ׇIj�R��]r�6��0�{C�*8Cazq+�s�vq������a�ꞑG�4���y���eֲ{��<���c�V��v>ī����+%0
��V�w%ǜ�x�5�4�Ml�"�K�4.�ZU����� ��N���B�/:'�+�wdD�+�	�{�D�D�1Yp�.x��ruV ���&�@ʘ���*7屵zYB�>����㵣��b!���-��k#ҙ���]�����Y_ 6��־R�D�]�a���u��fH��pC�!���5:���&�g��/�lI:Kc��Z�?�E��,�u@�\�ZQϔ��;�(}
�td��ƬZ"$��pC"��˜��&U3*`��%������m@h�$ו ���U?t�k���EV�$ ZL9H6�����(���ܺ�ɩ�d�t���6���ȱTfG}31$�Sw��M���ꡔ�����oE��"� ���0��X0�O��jI�^um�h+gՏh���1>iͺSZ?�K���6p��~�:FD�	����ס�0���6�D��:'�8��hw��� GTe/����St��sn{����@��U[әa�������)V����fK�a�8 -��ϙL%teNc�N+x�?X]�.����I)�$"Q������Z4Y��Ms�xG����nGo�@�鍶9��?����x^�n��`�;
�s�����.Xf�i~�9������%L���ޢ �8�K-�B�G:��9�\�%�O��x8��0�3��a��c�Cu6H��j�P�6½v��3����V}��l�\���Ӕ���}cZ+T����L�֍L��C����� ��#^geM���cq�PE|2��C8�"�v�-$��hKpuu��f3vԘj��nc�<0R�Ϋ�� �1�$����}�2�`SC�Yz�"���s������ͩ��vHK\;������Z�u�cE7�xt�3^Y����h,��o*B�-���R�����i�,�6�u8��@�@C�����ň�b��Z�6��(p��(ݣ��Q��L�Ç^���}�qH��-�l��U���w?��G}q��W�Њ�������ܸ%�� �VT�&�kC�5I?z����8��]��[~�H �Xڕ�l.�F�o�ey4������+T�X|MW�P�hc�e����,�65=����)����M��&Pwq�ԁLB|�J�%�W&��N�߅hI���Ǡfk���7�x|�ex/�CjF3�.#p�Y�`�l�D�&۷X�Q�0{T��Gwbx�M��q�<S�?��~b�(p�K!����20��(��a����Su�C����+����/����SDr�%d�֗�Q�(�Ҭ��(,���( U� @n�ڱqX"���ӄ^����H����f�8)/)�.X�����6\,�����7h�ڎp����t��n/��:��8g-�x[�XIԉ��G�:/�JP)S��rW���00Ï$�L�Jԫ�+Y����@ko��d]��`��`��4��۪rT�'�?����Xxj�pAe�L��yi�L	�F�٭�dJ�T>�祫��['1�Q�f'o�+ۇ�J�]�T�>�Ƞ�Ionn�x}���k���1漢�ã:�K�����#���t"�
�.�<�u������i�=�~`��HZ*���-�dt��ԁz]�f�?p1��u��A_��]}=��Z��T�ZXn�#"��"e�L�+b�Ec=��kPHDr(�%T3��ߘ��f�pX�>~�`E�aJm���k����H���p�.3`��g߲D�5���*�q�����_
�n� �H�Np!����:�,j ��8��R}�O�HF�,�.ˤ؆��������S��#�Ry�=V51u��:&�T��t�[��q�q'���
d`�����RPk/D�WԞ$�K�шrv$>xaw�����n��I��͒�vN�"Cn�0��BX�c��ŭ��8�Ay�1���-�<�D+�B��	�S����q.3j9�k�q=��T���B&���=�2�E��L���B�u�a���j��[Ή+D��1� ���V͉/�t+� އp*�]͉P��x�mS}V�,��NR�K��hп���P_J�;���/�ԏ!��� w�z��O�N�	����!|���pO�����w�S,�m@{���T�yQШ��f�o{�o:��8.���5\�=�˔�k�@U������o��k�����Q+����}�v�ѽƞ��ic/�i^���x����	KDA�Y��ͫ5ow�[_��e(��WCF�	������&D���/Cdô��l$1��2�>��Ehƒ8�,�Nk�o�)*��������޳Ai�ؼ�����y�c�m��|e��xH�V�9�@]=iL��H�R�����3�I^��r_������_�#DP�~���X|u�o�K��xD���K+=yO�z|OXf!ך���lH�����e��ˠ_�=���.^�@�𸊷F���܎�vm��0۬A�`�xte�<���
�pe�P:.F�e���p����C./)T{k��	�~���L�Cᡒ��9��S_QRD���54�:�S7�lh�?�]�ë[�����0��&��� ��_S!�&��߈���@m���i���R�{��d���H�M���ot�^���?l6816T��*�`@w*�uG��;�7�{�o
���0!��#ݛn@d���U���c'>Ee(T��+�&n9��FSI�/YL��۪d����� -�/`���M�����; ��P�G �d����|��w��\0?N�Ɍ����Ɛ��V���z��װ�e��y���lۀF�d�����Z0�{1V�ef5l��U���c鄷2z����m�e��tۖ9�L����[�#�����C���YE���Ύ��h��A�u�fuW{���`�[�3�-kș���ܵ��Qo@!��fȺ7b�V�D'�;
�͑�N��(a_��8ڼI+vM��x��j���Yo�:�ngA��)����hA��F��L#<�:9�z����ho���VV����3uq����'�\i����U�
�P��A��HB ��Z�F2[ʟr�m���"��4���cJ��vnC�W�);Y~X������50��*����c�&�`Е�c��h�j�z���Շ�-�����j~%�G�4R�4�AL�8��X�u�����8�b�x� �).�����*oz7���'&fZ=t�9�`���اf��\n��r���a�9��6�k��J(&W�g���[��t�s;&!�+q>�>�ێ�}�ި:x�(%)FR��r�&Ŷ��]"EL�b�*�����X�{]k{�h��a�78ux�~Y�J(]��c��A]��\�9�oB�����"BS���5;�!Fp���?zT���Z�Uk�|!ah,y�� ���N�՗>橜r~�-�����j���YH���Č�o��Y0f�}ݺ�'���E��X�����}���<q�򥸢��Ng�>�Cc�r`XW�:?p�K頬°��1�ʯ��jz�:N12���1�8#~�.���Ö:�e��2�VF�%��k��Ql�����	�9<���Y��!���:�LU����i�Iih��C4+6����e���͐�_5b�W���Il*+�\٥Q��s��/DH�)L��Q:�6w�}4�'R�
t�%��Vx��.���н��^^�B�i(�-��qKvn�y6�2W9o�Oo����9Cu��t�bX�_����3RF��]T�eM��p(�6od ��m�Qli���,ϛ�����. �`Ȩ� ��t�O1f�F��"�wǲ�6��d�օ�&���'���q�FR��N
��R̦�-�i@㛁�l�=�I9G��8��а"Z��6��I<��1�\SvC�m�+��0���)�/J���M7(o��Д��)U]ā�Z��������s~Yx^NڶAYqS$���J�
��s98鋏8�>=�Z�^�˸�$��Ƒ�?IJ��g�P.�P��n�1Q��[򜓟ߐp|9�r�wFU���3�M5�tE�n��c
�h��: �b\x�'v�����T��Zu3�#hZ�NY���\~�X�p����Zo2f�P�<Mt!�}h��	�	׃�1�#$[d��_n2���YG���*Up�܂��Z���:��i-��0RGm2\0X�d�-N�<cRg~:���R�{���%�^�{��)K$�RYR<���0俻�(�u�FG�{��r�RTO�{�z6�7�=�u��� ��QO������ya��En�0���������K:���aNӃ��9�UhʉҨ��0fK��o��|,��
�oy����f#1㝸jv��:Ʉ %�b����Vz�z9��b���(�K��������"��\q���&������U����5�]Af�rDD����#~��t	����	kgP�s�c`7!B��M�Q��'�r�U0Lx�l��r�X�(�Ѻ�GV���6�b���YݸU/�����	{=0��I��
�,�8$�_9�E{A�rƝy:ϓ5��"���X�dO�u�8im��k����;?`�98W�:=����	������9T��@��C5h�C��LAy}�ĲF�"k�(S�)!�Î����Ykoj�lx����A�,��^��[�"&'��H��TK�B�)w[�L6�7��s�췲MР�7��%��i@+���ܯ��7��F�*��9��MFjG�qz�od,��nu���GԂ:�x���q��L���|����I�|&x�r����������Vr�A�p5�NM�KVׄutl7	M
��0�\0r���(�b���	��R�q/�D�N�̣�8�>��:�NR�xVsG�R�Ė����^��WP 20]�Yy�X�K���֎܃���7��[��0���p�ļ�Q�k��6ںB�L|��ѝ��C��ͻ�P��ty���P*g��vN�Z⎐��i@���Z����A���RZ�c�ő�XW�ztJ3U=�V"5���J�����.}@Gd���-:~��IO �>�����%���D�e��T(� �Wy�A�&9V`�b�oI �a��V:Gվ�8A���j��+��)T�֧�S_n��x��đ�&��G[��!ഋ�D�����I!8�T�U^j��b��+���$�� g��+;�-��ZI?Y�[��v�Z��B��l�v
��!���ȾR᪩@<[yf�g<��Ղ�ܡ�(�i
��05�/Fb,���
8{�i�Jm���O�4�f�B9�Z�ۅA,B
q�m��PU^v t����+f�����tʘ �>�p�I��6�t<%B���������3T�L=<5?��;&Cr��������4��C
��t@0.N���/���=��H�bzu)��������3�I�N��q����8�J����5Ƌ_�
���6!������P�МΩ�J[7��D�)U�=����tME��$�
]>��Y�ưĪ��Pm�cΑ�S�븾8���1C��=:��6�-s��F��+#��f�e��gN@���-I�_�<���`*9m�����n���v�P/���yD�:�EY2��dK�U��Y!cA�)+Y��n�a%���Vre!O��@�A���"�zw�5�
��f ƊV?��~̋5����%�"�u0�dX��jtS&A��t+o�l���"��4J<�� �X��G�bbf�W�(L=Ex�<�5�|�	u�]F�?�ƺ�-�G2vu���[��k����Z��BH��i����t$�$�!�U���S��9�E�J��K3�]�^�4�^UZ�i���K���RT�,٩�f�3�[�KE#�T��iI�ֆ,�QM��Y�<�kSry�O��_mQ�f�����?#�e�%ޤ�ef��l�b�8ۘ�HC���th��!�g�� �k��r9v�_��#��T��ۂ�Y�c<(6�M���Ұ8�Ԁ�l��jL���ݱs�Y�H���0�k���x�jҚz%�1��y�Q]��k:{�[A��ތ��D�0n�	��|��P�0���d���Y���9Tv�=��z���k��6Y�у�����`�)5���R5䟨z��YG�e�F�X��p�FHcEͪ��۵]�u�-��6 L%��*���'y;0�e�m^��eߒh(��˫�2�l���׹j��6�0]1��.�4j�R�ݾu%Du��Γ��-�o�R���WlH�ڶ����e*�!{%�Y�"H����āKu��8g5�c9����pXH/�0�L:�5�+�A��|�y�i��nWA�`>�;�p��t2��:ł�*]����V��.���w4�����+��}��zo�$��R��y,0�@h�T��J �Gz�E�^���Lu��BE�:�Ռ�L���N�"�,T:c�����m���ߎ�xb���Ǭޖ[ÄP�P�)pv�d��[���zJ� �jxA��	XO�%���f�>>2����4�[8�R�޲�d�GX��?h�־a�U�`�{��~SA��p���?u�_��k����~ɏ���ƽt��8ݐ�&����K�s�C�&Ʈ��ٟ_(��E5��G��۹ߜB�2�j�N9� ��gm�p�	��s����a�E�q��ˏ��':��}�L�I|-����*Ë�E������m�
�Y����o��������z�ĚNo_A!�cr����k���d�A����X�wf�~«�ܜ���g�#���Gn�$�$��I+�ϒUB`�t�������囼�����78�	oޏ�1��Ǆ݀��^���w}�T:'����ޕE���Ͳ�����?%�O	颅F5��ٲ������<M��ExS�(�W����陵ZB'�]j��~@]#^����-u )�XA�=��9���\ ��8�5P�>����Y��=��k���@�\#A�y~���{>�9����8F�dJr��y�O6/.2��oҍťPN���;�=��ir�;o�85�j
2���cCtY�Jk��$�J��m4�`b�_?�_�@��0�[��`���r%<R!����Ш���C���A">���m��;)�_
��:1����;^��_X+�[sp�!ء�wWwe�<T�mn6#�(?Xq��'�����w�wR�� �Qp᚟�_��n��y7+����Vu�5ʳ�����:���G+����gd+^��,F 5<�0��R�"�/�^���aǒ�|� @F�F�p]`5�T���d�l����'��<n�$Y�g��wS�P��\R��o-�23�2�wꈥ�Wb�g�b���ӵ=������b%����`��&&���B���E=dE�JC�3�x�?�*���9_�0.Z�����<��o2e���St�3��|x��6�S9Dً�K�'f�5i[&M7wH���9]�q���$��m�l*o�{wRA�z�*�:ʪCj�;Xb��6>;M;�N�p���=`�oZ|�D���؀�[�o�TE��H��&gOL�V�qg�8v[@�vLg&�'��yh^)º�b�����sH�d�L4�ݗr�0����ݍ��!�0�ī�j��)�,x�؉#����� q���)��jJ�����߮��~3��oSסI���A4^2��{	��<����
f��M��!��{�t.Ԅʦ����
^�;V�,v�ӯ�%�뭞�.z����S7R���^h�\���&�w`
�{ۡ*��2c'k��IБ ����ZvS1�/D���%ň�1a�@��Md���*�<��-k�;;��&,�t�c�?������ñ�X3!Anһ��?�*�9�N:+aӜM=�&+���me]��Fr�g��W�i���j���նಲ��/O-�2#��'���8�׷Т��C�J"��a�>L>���B�ـ^� K��< ��`�&��s���E�u��&#vs�?*L�p�9P�|���u;��<h�3��9m
z$�tm)��r	�q�a�-�FpΑ@�nc��_�X"�B�!5��%|��L���C
⎌P���U9T��PG�?�@��R��(�0_�g�w,�0!&����Ԁ~#_q�b@�R��&�i�wG}��0=x�z�Ds10�>s¨z�ϫ�W�XxmP� %0�tT!���G	c�_���଺�V�a�t�R�W��4��^�s|*-�g�3�	��x�vߎ����m�>�7;�i���YVf)�DP�`������B=��t�"���!����'� �?������OP�f7o�Yu�=�M�7�G\w�zcQ��PJ��8F���"�}7�9�ֶK�S�	�~i�{8	�j��58��y�FݱC�&�N���u[�^6W"g�#�k��RD��Y��U� )��:���|�n�<%����	j����	��@{w�9����`�[��[�
����@ �[0�#��ܸ�d�?T)cٻ�w�Fz�x�wOh��ߕ�����4��������=ꮙBN���پZN 1I��}������D����wX}�G���	��H]��1{�2�!<��ba-�њߤi;n�������j���������6N҈잱B)��-�>��Xk��E��m!0������R�N��19 #K�Y����]������,'S!3�jֽ
�R��h�kn��S�M�!6"^����O9ff?�Nc�}��|�d9پ����w7��6�o� ��b�<�j֙�o6���]+zj
�����.���a�D�P`�	�z����{%[�`�,!,pݱ��Rr��V����m��Z!��%��ˁ�!�n�z�8�`/\C7���{MMmy$�6�\&K�u߂�;�WP�?ϱm�7�(�׷�Z�%n�X{����5}�}��QS�;K�"�	��O�
7		�T����N�V�^���\6��q$/��b�uL(xO~��?��ß���¥T#�K�|�x?����BO��I�c����+��Y5�HlFx}�3mߒZ���Jt�#b��%�x�d�kȾ�ʅ�R�ѳA{��s������&S]�b��VQǁ]&��V'g d�M�/�M�^��� _�&M��{os	��u�X�6ٚ�	pt�E_g1u�I�BJ&|�����1�Z��xv'�0P�BV�1E�aA?V��j��m��8������=�Pz�!�r<
�>ӗ�����>��t���k�Ґ�;��I�ڂ>q~`��j6�7�Pfn�u^��[��d�*�	���!�jT
"r�WqkW�l�MK�0f薽LyC%����	_��'%�وwo�m,)��?����&��)�2ǻ��ǖ�Դ���v<�M%�������q4�ʥ�R|�Y�����	�&�q#��V�jnB���d�3m̺@ֲ�*\�(X��J����.���H�*3;^�n��+
�	��c���vH+N� �����1N�yS'��[���y/=��	_�����dfXp��ږtW�+�~�m��O^'��j����?��7sGբf��� ¾]�Upcb����Q8 g� ��)�+Q�<jd�Vt�G���825NI@ߓ=F��	T�2���4uq�imn���WL�c�����y\L�S"��;�Ԛ�j�����W@E[�"�M��l�A��~\�MA�����ꂤ�KЊ�l�M���&_��8�`/�����v���V�pZ���V�H��y0�Z!81����I��{O)��kQVa@q	Eu,�pBZ0RB�]���2Վ����r�[��� ����8_�aڷ��(J����{C��v��ZB��X`C邗�{g7���T|3��kAT>5�\ ,_�ao3ѓ�TMX��0��Uf�ŘVC.N���}����v���Y�*��4rU��(
LUgMkoa|�/H[Z.2�-�W!�)��8b��*�zeLe�۔۾�l��Z�$Ve�p5DϾ��^5nḈ�py�� ��s�� 0lJ�c�Rnݼθ������j�4��ȷ8-�5/�bU�z����f�@�b��T¾�$�=3��7���[���9AYXO��O���{f�(���R5!����$��D'��>Ϡ�9]�?�̤��2���0/��mP�dp\P	���0����!Ԍs�[��GP5�/s�#w0μm��%�о�g�� ���z]n�ژ� "�(%E���i�3�`ѱ�6��ë��Y0),�|b(�¢{��>�Rr��Ɓ�:A�Su��N)�%�tS?�A�&�5I%*]����`~�*6-�x��\�yy�b��	�h�;#Qů��I�q?>q�Ǐ�8��3� U���Ei����	�6.���:f+� �]-!h%z�J�O�]	Pf i�>�4L�ݕ��Ց�0&D�:v�ajC���ޱ�E��V&R��	g8E3]x���>�$%��(����@�;�%ǝֳdz$��N�GA^֛�~��f�fUɿ�`YjPk�)��/�����r5P~��$�+Wٝ��=G���bI���D�q��|%��OU3݀�t��[h}���Q�uq�[��w���m��E����؍ �?D I�'93V\3b�G�4}���ݧ-���E�m�:��%��a�oy�,�@����C�L���у^a�#qnS�*��fr��Q ����vt��d���x���.P�#O�R}E	���Ǵ��]ď�v�4ϐ� �s�Y˞�x�	c?7����rLc�(�D�%0|�5 cR��w����{˔
	�m3۔P�;��Q����~��Z�O*��mbզ�����g��D��W�1$�~z^i(��D��J��f���v�;�	1*�-D��ţ
/$�?�o�T�M)�.�O�ؓ��	P��HTƋ�%�sp0��/>sp3����C���
�5v��q��r�;��e�;��jp������·'/Xy������5�r���u7=���%?��.���L�����K�����������t�u�O����:� FH�4<l��D��J�+��$`��ְَ��sZlRM��q���ʯΚ^~�rx�dׂ��"�~�kd麅����洬���dS���R=��t��zw][��sU��������X�\��"�8��¼���X���h2�&)�h��%�+��.\�Z�TL�=�{v:6&����^F[/;%J��+o+�GQxY�!��a.�,����&��σ�hHc��ك;2�]����Ջ��SȮ����� �_�ł�S/[�.�C./?ۃi߯�����&7[����1|:/�.ח���72�mv6l��
�,h�;^U�j]��Y���~�	F/�[�.�������S+M��lי��Y/�
B�J~髕-��Q�k�Q-�3�<�(�	(�fp6��2���O�o�(�4G�T�����O}���e��;���ۋg�*�]�zN�*x)��M'�h���;�E�S���9˹q�D���ĉ��|�t�`��ۋ��q����������A;�!"�n:lA�|��� �V�9�>EN��~x�z:�Y�2l9S�b�-�b�.��V�Ġ��F.�ްnt]'4@u<=��T�V�%H�9��j��ߔ�[ڝ�9(!ZaY`12nA�v2=�@%��}ѧһo1-�+a���x��q	q�c*	�;���Eڣ[G�y�!��������b�;�P���eߑ"�q끯�ޅ�7��6�,!͡���se��&:���fݪ��np�����_�ƾ��ӹ�<�LQ8\ݬuk8IvFm`-Gr�k�t��r��y�z�S٬G��jnݹ�Х��g�h���\�G.�j(yҕ��*�ŝ�4�D�R�b2�
m,��NwC#��C�[�=�	���D��H 4��S���j/;5�0�+�q��&^1CA�X%
�8-)��~i�
;6������+sl�#�Yn�{W�xlU��5��:Ґ�B��+���c�h��h�R�&�< �H�-���G�1�t����]ڃ�HCV/Ӎw:��ؖfm ��ia���{&���T�s 7���ө��S�a�f��gw<�A������[�ri�+�G`*�+��s��n��
>̣���iH���V�Bf�E�&q[	
����ik$-���r+�c������z:�w��͗��� ��S�.�A|� X��_��̜p�hT:�U�`�UkßT~&�_t����%��S�i��e��+�UO�[�m�"(�9W�B�j!�8�%��K��W�nH���;�
	]�+�����n����ž��3����r���o>�D�]GԶ}0e���Z�ɎX@5l���c��Z���, ��]����4���E/�>���^���}�Ć\|G����l�]��L\@����MPWb\�֜��B9��tV�ӆY�'�yI'}[=j�8Ys�v�2k�3���Y����J��F*�y=�#u�k�*��`�P�����R�uS3�X��f[A[�m�Y%��ŗ!m*}j^ʬ|��29j�:�J>�v�I���k�{��þ?�.Aj��5w�#X�k:���܋�������Z�7��S�yخ���բ�$��''}[&�UN Ũ��;�w_��in.J>� ����/)�=�邞��)���8���\���=�/�b�ޡiK����L��+z��p�g�gX\6~[I�O�:Tv��A(X�5�=�m��>K�Z]�KDΕnG��IV����8�"�٢�2n�b(u1����ڜ�FW��1Q4�B�W����S~2�CR�o�gvj~���1�*_�L�*�Cc� �\���]{����5`�H�w6�����ִD�֜�]'��Tr
�A�B��
��9��E�c�f�-��H<� ݀�c+J�#���a��t�$�c֞͞���/ӫ=u�s^͜`� u�q2w��64��ԯ�����k�N�r�Q�{�+�Rͮ�@�I�ze���|kW��4C�Z�V�C+���j�rŹ��|��Oݼq�XT쨣x�H�웈�h�0FF�{��-S��w�xl*V��6�%�y �f!D��
�)�f���dI1���Ԋ߆̲8DR��5!�!I_��
�K���Ў��#|&@m4,��x�X��De�C�%�Y�M���=x;@?	���~4�O�̞|�l���B~��[ �3�K��'�_�_�#��դ���&�;�4S[�la��n[���@��y�sW�<���	����#�w���{��csjX��_�B�Bw�.m�IA�6�щ^��©�Z��Q>}���h��$�����ʰ�@F�|1r&��]�!��Z�x����J�S�,Ise/�WX3�7��甥l�n!�9`��uIf@�ɫ<��.�P;�ג	�9��2���g�tD]�Q�����q-�J�'Ho�p�@���3��1;'ў�XB�4y�����,Z�@�x�\f�7Q���~�P�7l��ϋ~1f/�<G�NLcD~��ǒ +��"#o�� ���ΊY��ڧ$Q�f�>��\4�-���8=&���_��	�u%\J��[�ѣ�6p�]!K�#d�-Au��p�_+��pF4g�K�`�����f���C[t_�X��I�ˍRe��k(]r!�"y,�4�Bo���JI� !���N��`����p�[0������K����>]�v6��zH^�/:�~("���H�F^]O����C�3�F�7��v0�.���|UK���	ۤ�Pi[�k�R�+�&���H*���Q�\�Q�m�Pٸ�IX�,�$�p��_i}�q��Y2�l�HFu��-�%W�l�֛�N�c� PXyg�������sc���	�ص�C+�[����{RL�E����W�w7MV��Zs�X�!cf2�^>t�D���:r���
�ͪd_�y"4�kxa�L�L8�t����iV<U_4Ig� �oW����C�n�hG��]������%^����e���С��}��R����-�b���ݒ�kM�Wѿ������x�ζ�^� U�����4�mR�sߪ�X��t�t+ui�$��m�j2�Q�����g�DT��|	�j〔*�s�A_�ǎBġZtS�!R�m������_A6��J�Bl��:�p�W
��*N�g�6G��#139	���i�5H�)�j����]R^ ���0�
e7a�=0�8)��F҃��l�xĖ��o@�]�-K��TTkoC�fn���ݒ��}������讅��nY4�=�z�B�
\�>���S7�"t�`������R� _�>*h���Z4�k����D0�,����)̅�6�f��bS�s�C)K�,�e�4aCT��\s@Du̎a�B��2�dI�a]ܤ��F��X�}���'��WθEU���

A
�����Z(�i��e���H�!~-��R@�ƀ-�b[����@"�Z�)��\W���S�x�i�s�Ɨ4�U-1}�ׄ�;����B8e��Z�ܭ�1�=}�c�=ܪ�q����=�o&�P�(��\xB���s�4�^C��mv��V��i�%�����3��A�����-�cOImݏv�K�o�O�2R�� �\��6���Y�2�3S�7$�]�UyO&��s�d���i��gзd �D��j��s�� 8��ϟT��W<te�j=a����mo����>z��|����7�ih����J��{��\��Ų 0�j�w�r�f��;�o�i�'�����x�p� � :�� ��F5lA(D[.#S)�.����oa�<�A/&`a�CG�wU�U �x��R#dDB�r۝8H�*G(��VH�����n�&b��9vkO�OΣ�-P�6�'SO��a��\�ZY"by�[�u��N����J�ut��v��&G�V�l��`b.d�NX"�}���?;F-�k7�z.v
���+߮��+��������-��;
Bh(���7���7o
�>_�����
q��s0f���9�r�����'zp)Em��Kk{��9�]���Q���a��^�-&|��f<Q
��I��[�hU����`f���!����e����و�N��e�����EQ����}4n��V���N���fjg�_1�L��֗�21t�ܷ�ŀ��a�m�$i��x'�����A�؀l�.�@8W�],xz�ey��؆:��
�:Ϥ��S?�|�ʋ!x��ؐ'��;��Sc@����l���Ra:���Dn� i	��S�,�UУ�.�28b/r�RIWH�ﳀ��#�ws�"����t��eNʨ��FS\
�{�i�5�t�k���N6��f�D��`v�*� Gݯy=�@L	N-83����c-��ص��]k��R����vܬ�}~kW@�>�mi\/�-�`�gOf�����Fi~1q@6$a��J����|��N�ˋ �ҟ"A"��EȠ�,`#g���Bd���e��Wz��z��t'@�Ǌj��X�D�d��!�^q/j�7�!B�\%e�/���!_W�!�x���a�f�L�]Sĵ�"%E�'���\�}t��L'	yLs^O˺�h*�jb�S�v�GW�M���N���D8�?d5_qXta��6�Ć��9����N�鵲s/f�Q[��	$x��(��q,�ۤ�p�,B�$j$�r�߽}��nP��W�ߺ#�Ѻ���t�a~V-��}���i8��m�r8c �ƭ��Q���*l]���E"UH�����攤{��:7gߵ"f�4$�?۫9�����z}�o���-�$��c,�" o��7�_\ɣ��RI~�\V�P�lI<�8>>�K��|�-ㆾ%�Kd�S�d�0�e��P�3�uUJ�]!=�,��,?��|�{��!��Q����ta@t[S�|��s�s_��3�*t!d���T�
4�q�� ���jgZqM�Ж���G�����N�C;k\Q����đj�������{i�K,w���eM��j��x!�͹����jA"�
�h�\'�4A��W�������:K�bϝ��KK���s�Z��j,� 7���4|}�L��$��^���ӡgG�y����B)�i�I<݊�.�ɦ�	D�s,�j��r���~�*�i�G�[m��΃�.�� ��"�����P�����B
��Ѧ3����lh�	*��\���$A���a(XEܼ��5l�BB�flf`JX*��T���O��+�+HlѯwD��O��!����xy��Q�����1��Lj�=� ���=b���yγ��y-Ϭ�i�P4;��L��<���A��F��֕�Ȉiu4Z1j'�+T������g.�}�|�$OC��<grx��h�n:�2�/���b����逗rt����e�� ��k@<ͮ�uݷ��V�Z����MM4�����h������*��u����R�y�<�|�F�����N�a-/��Κ_�������X���tD:���KYy�D�$��������JO�������)0���%������*U$��kM�eJ��|������U<9�r��wo�ά5 �K܄��05�H��<c�7�鴘?3�3��"�F���"�Ӟ#�T�F�5$�19����]�r�E�q���I>�>;N5��9�/�P��F�U������xR;J}�p2?�e���4WX�i��T.	�i���em�6����<u:�:���Z���i��9���/�e2�āxMY���b�:��#���X�>+d�q���d�^��c�����ۀ�K��_&r��.�=�j-k��W=�S�w�ØC�1�*M���l!i�	����I�4V۪�����?m@��'���i��s7���38w���CN"3�&�l���j2S��Wf�0��Zu�$:
�x�/�R��Q�����(�h#�.)�?
�m�������FV�W����;�UYr�I,klZ
�s�?��B9V���/r?�$�a��N��Y۶�U0����5�7�A0��`]ĕŵ.�.~���`���1YM�]����Q�1�F�ּ��4<�d`Hו�Wc����Bgj���u
��[OAR�l� ���@]���9f_��Lg	s�����Ц)�ܸ���f3�(�t���s���<�s��T�����,\�G�w�.�TMK*�!��[��$�6��$|Rq�|�����N�����|I�O�T1ߡn*T�-�gREp6a����Y���Af7�K��D��p����$v"�)�[X�9_��#j�^?����Y�Y�qq�Մ�f�,��X�K����'�{DJ���n��l��}�+��;u�X��cZ6TǛ�M�7�Z�t:L�U�7`�T�H�q�˄ ˍ3:����&���8P�y��d�~�)��>q%�l;A*�������)���Z1I�0�u�YP� &e�c�$H��^�YE�0(����G��2��Uq���If"D\��Ѩס@u�L5�0����a=1DhQS���e"d+����mX*Ee(�O��w,��k;	 �光��mN���}5�����/��~��Im`���lW<�G�N��p�U؆��1�k9n���7H������q|��WB\���9���=������&Ş��@�g%H�v�����#IIr2�ӑ�1qFS@���P􉱆iOʟ���
���8�,AW���.$���>٨�~df���"�t���.�h�h�qn����}���$]u����l���6�JA0�\����k���B�a�����蒚�(�R���{2S#�J�;��¬ZK��e��O�c�.<Z��̂Ļiq���u�)�O�C9�xz�&6m�@��d��
�L��e^�0��@/`0|�N;�4?�v�����{Px����ѨJD��?�^B8V�����ԛ������ݜa�=9:�M(���h�'Lr ��p����]�~o�{���mm0���
�D\`y�6�*�����5�l;����<U�H��	 �i��m�~DevpA�S���^$�9Բ��z�6�M+���!� �¹�9@��Uo�y���iݰ^�M`}��y�tC�p�Ҙ'd2 ���3P��cU�xY��B`�<�����1 㔻P���Im�4f?e���:�Xe�ȴ��`T��=��B�c|���-��O}G ���l��5%)%C�A��z�K�����'��bY?��>����D;�Ӛi�����!�)b���tpvPT�f?� ��-f�$j\�{]��6'�4�ks�8��K��>�^�*W���_��j��>��=�J?���x	��?�i��]�N�%�w��iH�z���O.�0��=�Fӟ��Ԗ�Y}+����7��ƀE�#��r^��q�B��g2�������{�x�];X�6��	2W�m���J%�!�^i������N�R
�������N���J�o��'˶�~}��޷!��)�+Gj�T����Q�l�{��Θ褀\nsƈm;��є�e��ؗ�o("�L��'q	�\/l�!>.{6��Ȝ�;0����فu�T+Yg�{k�l������M�]�0��tX�)׿���&�F�{0�G�<��C�qhJ�N���m��S���|)ai�paa�6Y���<`�����BCԲ�3lY�Ժ\/}}���tE�3�W?}jτ-�����F/�����}�q[1kT��K�_����#������
�^���uFXU�бīUa��\����[�/����{�����RzL��@W{�k=����!�w�E]v˩�T�f��o,��-/�R	A[���Q���:�s��f���zʼ� r����MY�@���%���R�_�֐��9ݮ"}�kO�a��ה��F�ɖ��m{��|��|T���c�L��P��H��XdZ�'[2�W!�)Z�Ӵ��Gf�9��|���z/&T�6 �X�0�}�?(�g	�K��CH�X��5a�R07�!����J�9��g���4�pӎ2�$����5`T�`�Ùhs�A�E�S[`<�[ClLߵ�� ���w3tŮ
�&"{y�P�co�b���V��nU/i�C<�E�$�t4BWgB��`�mށl����]b��5�e�ˌ��\(1~���f-e_��:~��)p]1�|���^�(�m�Z��8�4�\_~�y���t���AQ�:�`��r���#� *Yl��T��ll?��-鄢S�4. %7_����ɱ�jM�z�)�l� ��S�!P�5m-_A�܆��:&�4�4gF�"�x��v��p�S�8�R�L���9�nt�<a�`8󤗍����b�p�9���� Q��4���`>�ƾ��&�������ZB�	b��W�Y�Hm���R8\HΒ�1>���U�-���%�2�@,�E��	���t���,y7�w�&�a!૯���xJ�9� �� R�Y˒��	����Vy*{	
,�oY��A%�:��:�i2�D��;�N�|�J�Ҥo���Q�w~�s�i�,6 ����Qp���}��-��+hi�@5}]���e��~�F�7L&V%����a
��M�t�x�~D�K��<���w=2��:���R����WA����b�<cݨކ$�������I�>��l�C��S�)
¦SbX�39PW��ޓ��&Ȁ~�
}߻=��0�;>/��6d*4b4nʽ�;�,��ce�tu��I Er��F��%�n�"�|$H����/W`��"�s~�pղ��YI�!{��B�F�EǲI�R#��%tW�T�ը�����0?��hm���Y��E�H���W���ho���5n�4�<�Tc�]���WP�w�^�����_&Яш_�����Y�Q���5���0=f�fN�7hySHNoW=q hx��d�gD�5���/u���>@�����=`p��UE.����i�H�"����[��]����Eо,d����[J|����(B��&�I����{�+����̚Eu��N�;9cKRN��t�O�	�����{F�+�~���q_���#�82P�������~��{���Z^g�i�a!v�Ȟ�{nL:�c	Ǩ�ӄA��!�����˼l�x�Kv�Y��T�E�-憊�e�'*��v��;������R��v��>�����we���^P~�c�>&�M�N�/]� ��ʺ@恠?j1ֆ/o�=�dma�G�)�-�--A�x��gp�v�=%�Ji�W��Dz4 �K�2�@��0�4y��6ҭ)��:��=��2%�����;O�3�5a�'�=WR����Q�ԣ���j��	6i��V#�ρPqT����I��B�Y�t���$�5Y�ؒ+ֵ�P��UW���r����>�T q�Ӹ �g;�E�GC;*��	o ���0��Sp�ڌ)0ಪO1+���˩�Z��w��n�b>x�t��Њ����.���늜ԽXDݨ/������i��z��P>� �����Wf�|wӅ54�}Sv��{��j��M��gߧ��C�S����
PH${ �o��C���m��U~M:�QfRY��2B�}¦��u��iv�Ի�b{��4FQѽU������ ��1 N�c�E9���Ui�����m?NBF{7gm�-$PZ��|�5�]�7W�����L1C�F�߭���K�{>�i����r0�P��*��S�ݺ��gc�ޜ��l��"���8	l�v-CީS�k�1��+깱�L�tc�V�:0J1�2�Ӹ����Fwr�K��[��.cεzt��+O�Ypo�K� )����u~yc�瓵��V�FA�hv�������p�0.!L�K��P1K%M���c��Z��(���3?�`l�|�!�;:���z`���W�Q*~�B��J�t�=]!:&�@�Ф8�Q�?-c$���!�F�EN<>��!%M����V?��P��Luw:t7���=�Bhy��	�q����g��Ta� �Z�ey/&C�v����g����]p�����������{�C���Ys��Xz=U:~�V�������j����rhsp-�@T��C�ٮ�U�$�$*�v�$��$3z��["	�\�wj2�����x�T��|�ϟܟ�>�g�zQ�S��yswUnmk�ݐ���j�y���Q<�����/�#.�6�ߦ�t���$��;��s�X�a�L\+�1��җ�g3o�5�t츓[%Aui��)�CE������D�59���X�C-BmBz��\��ł� `����̚oN{�^� ^5!�7�c�����W�5o��<k�m�i9�����gˋ�2�Y�)���B��E��i*���ﱦ�K�敚�"�v.�+��ǆ�m���I���q�"[E&��5��u��_W?}�����-�?wӴ%<��E:R�n��ɐ�x�|����Pk��5+2g�I��{	w��B�ż��c�зӁuv��~89�(����>��Smmi�)�?�ڞ!k�R	�K(���l���,�1���t�ܫ�:���$\� W�r)�aYk�	���Q�mI��m��ٶ�_�O) ��IgD��+��dK��s%��=Lٗ�/���1L6I��
s����f�w�v
͚�s�4�f��f��~<�0�E<0ݿK2"!� ���aʴ�?�
g��L�+�����J���I�`U���3Z��#ߊ1�A�bN��G��I�g�d1!���B����U���y+��x��[ ��/K��������)��d�{�%qY7�o��%y�T�+:������;�K-�bu��D٢ڧ�����m)�	r��S��� ��U�(mؘ`8M�b5��y!�շf�zVx�a���,�ERIX$�B�.�]E��5y�����LE��qbͳ&�0���&k�aH��f:�ZJ���~(��Ț�*czN� ɶ�\��=��9�Y��U�����,�Gv�>��w�=�ڋ���[�`*F1pӛ D������k�A#&d�>�����i��r���~�J�Ҩ���8��Yg�}q�:��4�!iI�T�<�f�2;^A�i��[ο{�aPK��D��"N>֡����L3�9If	�F�i��,��2 p_ Jq:�Qc�; �E���);)X4c�x2k��ɹ���:����|�{����[F3�]�L(K���?.ޣ�;� ��	��~7!�P���G$O��c�U��T���� �21JD����)�l3����Z]$��޲�Qè�����oP�}����t�G�<(4�j�@�ff�/WM���#+˯�b�"@�{U�7Ϸ0�G�F� 蚴�Ah�ߓs�Zf���J�!V�!�˱��WR��'m��Q��N!�͋s��b;���:�B�*҆y�8
�@x�����4��s�9����O=y�rܪ��Q���������z�yp��\!��SR�I�M����l�F� L��r�G���y{�t�qA|�i��D�A�?fi�#5P4�`��~�>�]cv^8ۑ[�՞���jF�`G���"�HX��d!DP(�?�Bæ����w��;��^*D�ρ��,����r�x��px�'�,L�o8V�����2��{��7!���Lx���#[`�KȮ[�il-g{��͉o)J+��M�aL�������屏���q�ۋ��.=Va�6[-����KD�-��<��Ӓ����%��tJ�������@X�@qfP�Cz��Y}G��8��#f$l~�1:���٠ݫb5�y�⦴	���#zOg�d&�7��%Z�xl~!icc$��V��p�`Z����H1ߊd�f	1]�`��ƪ�A�7��q׫rυ�����z����d�u�o'�!�E�q�!"�H<K����Ʒp��Zgz.��f=�"y� %�؝�i�VaN5#g�Y�bva�[�������E�uĂe15vp�3��6�ت�WyÏ�Y��^SK��q��<������U�����+틺�߄��yS���Ix�-x����!���d|4����(�@�в�=�o�uxV/[�I�����<
=����?]@��jy����J5SNnlfU+�*>sB��ٕs�ҡ�3+'���A��u5݄��L���_�����͋�$b��#���)勔>�5�v�=`�����F��x��oޏ���_���>���X!)�z��̌�>��r���)��c�Y�f���?�*��ڮ�	s|D��עOX ��gz,g��eD*,��Oi4o]���/�Ň�r���v_"]8�\L�����7�EF�M�kȱc�[��;�\"��iVO0��=���b�'�G�IFܣ�<��R���a�~�%p�z_|���(����׌���RB¨ѷpJT�B<�]��e|\�Zd�v������C1
5��l?�e��D�_�RP7b`�����@X'C=���%U�,$��h��i��:���;=
T��+<���6#�Jk�~�&�����Z�a�z�3{ְ,�w��6�v�-��5���D�:��y#��x(���;a�'R��|l�;,~Dyd��:��G-�4!*O�s)H���?$q�<��#@]� \m�A��)����V�bq�<|,�7#X�w���ܾ��K0�o�~��p��>l,�\-�8G�4��Eq��Ό�贊.�/��ҫ����d���Fvh<¡�,����5�6Т�J�#��
-xb� 0�;G�E����eo��	 Y\�l��zS��0�[�3���;���5pZ�u��_b����V��H�HUD�!�U�:y���
>R7��w�c�2�(A#�Ë'=/�yn�����B��օ��,�j�5��H���p���B�{4˃�&i:�����5�m�M�]��������]�U姙opω�U5 m��Yћ�5\�;HH�ŝ.��&eI���I���=�&c
�4ʝ��d�Xְ���5���f�0� �;�|��ʍ�&̖�Wrl��AIa��������2+�758m@�c=�a�9��I���h����$"�?�Px���@��%��:]!0X<�WT��X�p^��G\���-1�e�檉^�dSĴ`�8R�,R�;�Fְ����Lc�-��<��o�X�$F"줼ov�f��1�̨�<�"GBS�3_)�߄��vKH�'স+K�%�+M��x�h��$�x����ۮ+l$���@�2�Q�b���rN}��iE��z1�@bJ3�ӧ�y�8�W�Z��OO]9E&G���C�zX�f�Fj�s	Ǽ�Q͜MK5��>�#�y�8*����R.�"�������s <n[��HSre3��K����m�/��ɥ�du���,���+��M�|]�%'u�6b��vƮ��*N���P�5=�*�?�|���
|0 �+!�!!���@�>޴5�jph2J5��x��e�lEc�7⯏��G�G,�eD�Q���D�ӳ�X&F���2���wE��(]���'�����tM������/����ǘ8Ń\=4��)��v���߳�YsB�SQ�%����@�a����k4����r����o�l�ԕ��ա�w�
����I����6dI�E*qz��*�D
.�g�93%��2�t���
����cN�r�饲�,&�x*�+���}��ÎvqEb�d ڄ�{�h���h|h�>%l۫D �mRVP#������U�92�ei�N1yU�/��A��P��|EM�
5�V�FT;���*"ֶтM�PtV�FiT>Nx����CrՎ��(()����kw�N�xF%�&nQ�����j�Qo5��B?��?��ť��jZ�pN��cpJ� !_[w]����HY�q5�X���������4�Y�����Z[4WJ�p˩�B�����a_�4U����?h��$�,2+����CY���1T�3�+��˹�JXo��^%nkɑʎ�(���0Y*	o�+��^,)�w�oGq��(ᇮ(f�%�T��.�Y�ǔ68�|L����x�<��?����ځ�]�Q&LR#�e�(� Grx0�fĭ�������;`y� ����Z�M�E��L1�[����YU?pM��S��w����R� k"^�2��s;�j���j���A(g_:�nۻ��J �����E����f&�x�����/���/���
(������>M��W2W/N/,}����9ݿ�S��7K�z�M���6�tv�1L�cU8�"�D�U�
���"Tݰ���/l��~�v7��K���x3P!-Шw��EG1U�K�nĩ?��;,xMw�sHW������V|c�z"vw��[k|�O~-�e�~�b{_\̖Wv��Xf�ia`$�_�}!�����B:-�p�p�%�ԙwɀU�}G(	(���EE�d�ٽ��1�L ���{ߝXC��?�%lS/S�����kmC�����n�ݼ[_�8(���e�(�ĞRE~7մCR8��,��}lK�Xɏ���M���H�ÌQA���i�S�^�O��/��'��2:^�� ���}�P�7#�SUMm���qĆE����
N���z�㙾ݚ�aF���J~��'����^��WB�YL5��������,IR�h|9��AZF���G%U\�n;@������#�����-��A���p��
��I̎�5�}��Bx�rR��_¨���� v��k�Zԥ��<�iE?Ӗ�9�k�E�����^��szW��j���Y�t������/�y2q���բ�Z�J��΢ṟlk'���dCh�UZ�A^�MK�NDZ����&�Gqcd��t�W��L_B�]jG�un�����/>�aW7���i"���X��?�Vn�_�\ǚ�;d����۶�k[��h�g}J�%ɐ�#���)R�Em�����1��Y���6�(�� ��^���7��?�u� *V����H�@�s<-���84���p/��F��.����Mb���bq�D�tqB�{#�AYin���i[! ��ƁD|I�w,���`f�� �q���
wa�Io�&i�/���\$(Rԣy��-=-�l�l�����a�S�W�j���{��TÒC��o�dG�~d�c��!��I%��rJT�s^���������
pl�4�tZ����'DlzO��d.�q]�(0�P@VA�& �7ϩ�G}0�c�7�W�p|1v���Y�<CiG���`�]u��4�0�w���G��I����g�+"����!'����K�k,��e�c=��ڊ��g���7�E8lE�b�Vv��l�����X���L�G5\���L��k6�`��t��!������]�ߋ�v }��ܼ�oJ�>i#+�q�r��MÜ�jMk�X���o���W<���"���-�%.��n����_?��x�Ls?�+�<���-�#�2j�G;eH���7��r�1���9����u3��dӟ���!�;5k�ԕ+Rp��o�e�
ӥ��Ҝ����7�W�L�Ѻ.�(���`��YM�C�j9�oc�6/*���9�%CT�
�"Ru؈x(���!����uħۨ~<�I�ʌ-r�EJ	����TPH;#]K�8�z�(�5~�n��Qk"��=�{�Ef���Tf,��v_t�o"Ht����<�Ȟ<%�>�l�tm���:�9���IpǛ�GN�{�"�f�I��?4�UE����k�Ѹف�o�a���z�qyg���=Q3l��dd�(\v�r�A���Z�믆r���Ƒ�	c�����x�����u.K��*��'��Mt0�_NЎ_H5��aP��Y�0�"�&ъ�LnV�A+P9T)/�C+^P�yV��`/��g��q8(c5�4�"4gH���G��)lJ����f��#ȁ��V�13��r�G�ʉ+AO%d�6���	���.i���]�Rɏpd����w�]"y��2�q�'����k/kCF����*�z��2��T�fm���7���+�{�Pc���k���h��Vʺn�6�CsQ�|DS�$
R�G��3f�� �PBh�T2�zb
���R�ވ�E8�=�W*D�>q�̗x��^�hV�!��oԜ��*v�k_�S�==��#`\�ND+�K�Ŷ����HP�>�Yt�~ž��������09�#y�rb��d?5�ExZDo�^��fL�?e���ba�xN!s@]b#!�C�=�x�l�������g2����6��́������:���5�W8_B�3��$�� �:�1�Q�����lv�ے�8��먟&��=��G���S4��Xy<�F�����/�6��1�Ո��Wy�ɸ+H� �~�s���'7����jv2?��GZ	3���0+�ג���B���d�}l��J[
^,�I!S��x�����PhBm�xY^&���H���OXj�:G�vC��������Xa�
G��C#y��L���e���y��
�� \�u��c��1F����`ʗ��39W_��+=njJ��?�����,?���F*�4]Db�̌7Lw)�Њ�!Qم� ��n�N��j���u�Ջ��,g,]�=��b��NOAN��t,><���T����OEiw"W	�!T���@��5<�	D��!�?��#K6j��m(Y��W!������a��n�1��@��=���#\P.�o֔�����^���>4?��&oѕIZ�n��\7	!0�U��^S���O�	��ʘ�r1��j���E��5����Bࡠ��ggb�$e��*e��[Fv�ۓU!qLHZ�a�q�Ja��G��(�Ӟ�����T�#��gPR?^õ�{1Yq���,�NU��?�d4-����R.#&���f�C�9֮��to79[�;U���%`$=�ܬy�l��e��j�Q��DD�H1��lĚ��X���~~�S���2��pq=�)���H��&آ�z`F�C�y=�V�7�j�c�P_{����������zr�Qxi9b����h�`���_a���Vm`L5
h�#�ջ��Y��g����2Q3�i'�Gt
��[��}?8j|K��'���J����b������M9u��w��i�( >�K�ȇ�t�A*���J�h�D� %o,r��^&���ĀRW�D�n�>�M�D�T��Ϗ�ٵ[�p���= �*k�xE�qu�������H�ܕ��f;�$��z�jBL&�m���&��=fO�:����y����Ϋ��v"��`���.UXR��+Q`k୨s`n�&�ΫI4��g��J��!O��oHE�ߨ�(��p���c/�LE�����C#�YDL�`�UL	�㩇w�3�A�� @if-΢��{;��Bf#B�(l�t@aA�mD�'h:imL߃��"���|�GLh��S���v�����~C�r��u��!�������HRK�C}�����_SoKr%	(T	`<�Rw~.�yl:��� �>�o(7�5>0�OP0����d�b�Z��w#�fb
e᪚����;Hg�8�x�[_Yq����� �S�ΓPp�N��.pbAҗ\N]���ĒQY���f}��TE�G���uj�Y��.��J�f��k����kD��"�:a��GPh�ԫ*O��y'(w4���ݮ�l@e�������TR2�:8�i���BgԹPc=*��L��N��	��=�H��96�&�F�/�l��e��!R��S� ��K��Dz2BǑ���%�đ��v
�5B��k�Y܆�>]p���^kۑl������L�1��aαQ�N�TD��?nV�>�]���',�U�g��t����,k�@Pm��Aݘ��NY��~hn	��.-R%��X|�������ݡ�k=�5 Rs6`�ٗճ��Эo?U��O��>+n7���8"عB\����3��i)L����t��SN��4_C@;ĝ'p��@31��Y�I��@�[�vs0�jv/��A�֡rMw�<Ie	?+F����7���l��	w��Ɛghu+pj�U��̕�b0h��r����FX���-�'�4�/0�ҥ�SE45�Em�^L��:�]�B�;e͸|�����E�4kZ�]%V��&G�Xa.��×��Ce��6��������¸���\dr)�u�û/Gf�t��ѓ�/�9At���0�W��ࢁ��T�z�}�I�&��ނ�S�����J���*���^8.4C����X�Ӻȸw�F0���Y�˺�9	��B�>%<GM���A��XLw�aŒ��b��ã8�I�3��׼觡�[8(�?�+���| �� K����xZB�0#�[)5|�{�b��P@�U��*^uK����X~DM��'�;�����)1�&q�f�eBN��J2^0�*�#���T�P-Q��dkG�1���P���`���#Ŀk���M̦�c��/���A�?�� �׍��~��.�'�R��y@ :/�`q��~���2��z3�w���DK$u�zq�,�
���	H��K�~]���3p�zr�/�W�U�����V<
��`�|)� �"b�9��M��*������g�f� �YD4�2�6�5�k.BP��i�\0��[;t�3Ӟc�_�w�p�sRn�îx�	�V��l��E�˚��p��iۿ3�'��ds����H������$��mx>�j�Ň���п]�SRή$��y#Re�$�zZr8��]@)��x�Y�i���3�4?f�gD�����d(5�g�ƿ;��ˉ�z��t�������ʸlc�*l*H���dE�Y!�B�DT+�m��Y�kS�Ӧ�l6B�6O���S��A!�rÓ;Ny��}��L��г;=�?��Z֐p�H���E>���t-�pv���~�����q=f��H.��}��a;Y��>�A�� Q�"u�>Rq�{�eg�7x��L :)ѱP
Š`�C6���3�D�/�����]ܩPmƖ
��#���VI"��ѫ��Ai�p٣����5{Ց�]Ee��kc��v%[��H{ܓp��ڑ�
�|�7�
��{";N��iY#��x�0؆I ﻏ�@���+�I]M�_PR�y^�.��OK�/�8�AN@W�Y���jw�ˇ���"�xǐ�~��T��-K
�nvJ�;�Q��7��$Q�TM��r
��-`@B?���T����Z��TE ��ϝm�ߔ��E}'�����e�.KL��"��% �G:�3mI��9ǁ���2��B,�Q�+����� ��@�S��5�v隽���g��ڽG��:��ң��M�Pز+K�-�&1b����DK3W�,؝��X�'�?XeǶÝ���u����������Ϲ�>p����p45��!)$!{y����<؇@�R�f��52�q��8����H��Q}Lf�8��Y���i$�,�����L�^��:�!���L������ْldɪtE�?��&��X((�Q �t_�����S�5)��Ô��SO=�<s		yU�n-��n�Lo][���^�`��p���4_Hڿ)�ꌢ>)Ƈ�.xG�Y(�0�x��5�]�/I����C�����)|�)Y`���\ȴa1L����T�-ѽ)n�${�愒Z�;:��V&�G4����vd��i�מ2t�Jƽ�-��JڛX�:�I����h8��M�����Q ��ҨEw=�@ F$��O���$� ]�j2����� |��h�O��&�[������f���5\[�\�l>1��޶�S�/�3�l�+���.Y�f7��w��h���Np�u�L��i�O,�P�E����?�	0����a�o(׽h�Qm�۝���]%^Ug�M����s���$��d�קH\A����%�9�$��/�T�=��<� �2:���*̩�yӇ1������O�@�w.�׋M�\����ᚥ���1�o���G���;�h98����9J�^N�<F��L��V��~ʔ�R�yo{}1*��.�"܅R"�$IS�t.�#BE �E����zݾ����p�?�4ZjGB��BC�80[6�Vغxט;���y�D�u�����L�S��� ۖ+��H���\�mbC�X6�� 	+���w
&@�z`���{��"K֭%���21���f�&���d��<.{�GASt��Y}zFM����Z|$�|+���i$:5�>��g
�I�RB¢ɞ�j��;�rZq �cB�־G�^tL'���&ao��g����s.��䢽�N�;�m��8���:�`�e�VI5Q관K�J�YM�:��x�BU�W���ʐ*��K���Z����E��kO�q[/J�q���vzi���W��Y����^s��:4��B�"8���"���i�?q�6�2�v�e-���&Ed�
���=�
_]�к᲋�cG�/r�:H�3���ʓ7!����ך���(M�x��pc�G�ɬ��}*���y��\S�,Q'5e�6���mH�VXy�#��lb&��6������L
�<�<���d�u�c����-Q�`QZ��5�������2��\?͓2g��P/��_�h�FId��T���e������Ў)���
2,-�wҩ�n�)R@��F������φ䄍�ha"�#4�HT�G�l���M�]z�%��aj9(-�^���3#�i~��w"O�'e�y�m�·fJ�i��D����y'�w��%"ecQq��:�QRPΓ���)C뿛�*^��s^��Ysȅ,希~�n�.�� SM�xcS����&��kӠ;����u�u=+rz�WT�UA5_�w���(YP��^!�֓@����&���$j���f��a�֜s� ��!��ʛ�R:�M9eRX-�,1	�!���.��Xp�*Y�87�I(`�Tq�D�$�/��503"��:i�.'�|��*J�*L;Aˢ
��e`HH��yܨW��e���[�x4lw�=pl��r	&/֯��4�k���S�}���)mta�$n�!H�]}������P��F�x�o#Ĥ��C?�]'�A��3�B�Z!j��T�S��D�pW�o���q�C�xf�y*���+ʺ��0z�B��3`�ʔ�����
��U�>�ɠ�p'~|����RH킩�/�XsA�Qk�+���HqX6�h� b���M:bnܳ�#P��Gw���8���R�r.���:ۨ�w�Gzžy�'�>�O_�#
�� 8&��V�J���::Q��k� àw&z{��Č}�����#W'4�	
��m�5Ξ�+U�� k�Mߖ�qV_0�0	�ב85z�>�(WPq���%�)]�
���J���j�H�hg�Z��`�a��33b2:b�c�խ�N}����z2$���wk��N�!ڿ.��pf�q]�Px�ά����n���
ٍ��f=P��d�c���\���[�k��;��BTy��{�����U]�G��*������!�ޅnc9CL
�}2�O��F��G�9�#�HKt0L�����؁�[�>H@7�.x^� ﻗ�����E��X��e=�8 ���z�C�s���C�~�7��?�?���eF�ʽw��lDy�Jh��a���ԃ{�BE�н&=9��"wcF��Rׁ}.�[��M�7#'#���@�Q����'-"略�\�,&�|Z�n����5~�2M��7�9��l�5�
ܫOz`#�4n���q�������;�ԍ��[IW�p�J������x;�'=c]�]�[�����݄Hn2��ٲ)c(ƃ���5��܅�E�� �}��$�$V�57M2"����G� �F=\�{Қ�h��L�E�(ؓ+n�2���j�3PQ쩏g�AU��pZΟ��kӯ�B�����T��r�-\���a#�y���c�}�������{�Lҟ���Eư��a�9PK��=AJ�j{[�r��r;P%یcǐ�����{�� ^�«㪔��.=����9PLzK[4��t!����8�jT83 $�����XG�ᦐ�~|��Q�څ!���u196�.�����Q�ë�B����^f��G4����MW���E���O[�V��w�������k����oZD��[��Ea�23���l�Pg%�0	>򬷀���OT�����������dj?��h@�W�ܰ"�N��+�\Y�����F.u����{�=�����J�0z]K=.E��Z���ƫN;�LJ��N��E*��<hŒ�6,���k�>ENK�-0_^E�;��A�:e�ޑ[그����W�h��\�T��$rM����q��FG�u�c�!HC|���U��j���/�h�g�zI���x̫D���b��u璆�#�RK�c�����]����j# n�藽;�:"ƻ��o��@f	��>�na��M:��A���Hhb֑Gµ��Xt�?e>�lBFC^�;J�8|"z��8�e�����'�z�R�zE�ʕ��0p�9��1fz:8�^
��C�W7@�כ����LX���F�"�M��XZf�jL�GI���E��:Ӗ�qG��	g�ky��$�C����
~~tK#*E�,E�H��R��tHP:�`|�Ɍ�*����#8�kP�v��j� ��7,������۩u�z��;�nj8Ď�#�mň�!���6(��4�ۧ^����b�]nJ\�;ʺt�hãE�'
�Q�8/��5}�4<	�]�|�r����s��[C�����,ӿ���QC��7Fd0E��w8������/���ga�>���D|>?��G",��AF���\��[I���S��@T�zQ�_&��x-rw�bX�g�@9�|4�I���4mS������>[����zj�b~;��ս�T�1N����PnD�?(���}�����C�Hӓ�p���Ff�����OT[6Q�ړ�������ˇi��l���9p���@�]�9hA�Fj��]d^5���aS�,��Ҙ뭡�>`�
E�� � d�? �*n~Z�V1;�	�����M^G|%8r�Y��x���e�ҙ�3	ְ��J/DR�V�\��,�6�B�^yGXFI����ݰnל7���"�Hk�z5�r�;ݻ�j�v���ni�\8� =d��?���2��[�?�K��b�$���C0��#�^�p���ů����i����w���cf������kJ:�Y� nwE�7�_״Tc�4C~h�w�J~�v*�]���>� 
��ޙ���k�KQ����:0�	��q��bL�ix�<��C5�J(�d��z��a��?%Rp�?�3vT����1��.��Z��<�?��K���l[Ž^�W�ىI�S�1�e�Mo�ɿV�bQ�蔏0�
��u�Iʦ���[=��E�5|�I<�?��Y�*�Q�L��k@����*,J: Uݩ�[`��(i�z*��w+��4�?9�,�-����+B�����&�!)���-��-s�w���ܐ��b�,.�,'�u�u�ƩI	��S�@z6�o�[�B�iz��R.�ܳ�\7����93:��r��tXp�;!6\����"�+���L��0g:ȴ�8��Н�N8�����KE���	����Y�Ն��T� `Y����j�Y��9��ޙ�@�8��KW>)�Aps�JeW���z)�|����´��8���nc
�9���t��T�y,��������K��F�Q�R�_�+����y��h:�#NHr��x9�Ǒ�!!��T��=����6��a=�D����\<�9ɕ	�
�?!�䕭x�A�leLrVJ���4�H�c�!�v��r��P�9�!��/vtF�P�JQ���j�-�3�+b[�e�ጦ���}�#U%Zj�b���A`�,&�QWPT�r�h�S�Êt`��Ǎ�� *!�`*�?_e� ����b��t��]��Ztt�M��K���F0���OsO�~�/���L<I��YJ���3c���}֥E:�T} 8K� �)C��x�^>�&$b�ʹ�C�+����T��I�M#�������)��Y�	�mE
M�ۿH`�,�m]e;��`d8�w�L����0�M���h���Ej�im/m�$/�fЅnl�/e~	�oX,��)�"?#A��qZ`$C]|F*x�J86�<�O`9��R�]|8)*kO�0��AN<��UR^�[=�#�������?����86\L��]����+�x!:��$�yY�b���:A���s������ 1~�q:P�)�V�x9�t$	d�R�%�
=�XL���𶖹�]�~�/����$ �d���N�G�;���,�/ň N��s�[�kx��x~T�7c�P�Z�^˯	:ǣ#���Ž�l��뢚8/zuCpw}y���q���Sup��c�&���o�?�Rs�"��/ul��),�]8L��D5��F��F�r�ޘ���>@V_>���v���n׆�u�Q�$�b��0�#K��&+��ۨé�<׏��(�u�;����R�:�h��W���t��e>Vq�ĥ
�K�ˑ��ɴGOɶ�mFX�d��Гہo&?}�C�Xx���ȓ�nm5w�wa�����[Ԃꫨ�"��ڛl����\&M�GC�
���{�-�~��}���'X��d��O�)B�꘥Q���$x��#`���qy�5)𛝯��kF3��)��74��RB�}��+E�!i9��
"�3?>���1"��Wo�[��C[�?
���_�7� n���������Y{� �I���˔��9��'XH��!ӊW}������o�3A@���Qb۵�v�"� PaM4	�u����?n���@73���BU�d��֕�̓��s��E��������V?O(8���a�I6��E���mgg������"���	��uWA6n�4�bYZ)�`� �@:��9Q�1n�J�6�eQS�y�N��zqU�C��z
p��=ŏ��9�m�x��4z8�F�W;fS?����'G��+��_��]�p9⪬}W	ٞ_�N�zrS9�����~�n��
�IX��A�O;����Ɨuk�|���b�,c<J�N�lǵ�"���6�I�����$k� $�T�y�پ�4HY?j��jl��0����s~6�T���C�C�l9=��7���m �`��w��Wdy'8���>��5���������zCl�q���~��	�7�} ���/�K��/���$==#���X���Pt�&�gSX�?Z�$���n��D��xpD��N����o�9�Z��.���1�o=z��m;���(�Ь�I~�E�꧀|�}��d[����So͘+R�9P3����M�!̊����^�E_��qx��<y8�x��Y)F7�p��%������&�����C����Z�S��Q���x/IZ��S'vy>������������Kh<�C]R3�8	R"�dh���ŉxgE�-�n���������)�4+��sܨ��*dR�P5<{9Y�ՠ���q��e�𝆑�R#E��{ K1�1���Tg��jl�1z�q J�D:���R�~]��%\�"5�ꮅrZ$V�E�(�W]2�P����^�:�b0H���#�����{�@ѓ�r���h�F��?٘�Db�n7��{kX�v��w�j6(%��������jHo�s��M0��5d�_�����@*�E#8���(ON��"�C%ta���=��cj�8b�S;��
rf�V0���@9��+t����Ջ�YB<{��j��C�[����V��mH��{qcf��%��2��j����L�$�@�ɸt��ju���1���H��'�?o�Tz��S�8V,�8fXS�AG�?����*.���� �����+�I�Q;a3HW�����{�Uе�v;"��Q`[�8?�t:fyR�'��@�E<Q�x��+r'w�aD��!C�a��+���΍-*$�A�=8�שp�p������?��%1Fè8�=�m��o�0bP0m[�blbV�)�ÄZ�^,ﭖ	5U���ԅ{��u��5bf�+�<ȭ@�ܔB:�Kߖـo���6�@�A,�~�]T��{|��{�J�"ƤI�v]����xqya�i�*�M�JŁN����4N�#�}�/E�LF8�c�z��dӧ6L,����hvcP�QUc�D�̿	���oH^�z=U,Rg�抶n��Іj���k=�U��Yh��k
�nDc��~N�Wy�0m}�a��~�E�ݱ\�U2�*�{^�%$q��;.�*9��3]�)���z5���j"qr]/���1��g7���hwPG���fX�LέM�A�e�ҁ�şz�dʓf�O��Y?�L�l��UZY��5�xkpx&�#٩,S�ih��;��6����g�>�L5F`-�PU���F�pᓃ�������/���1��<�/�g�i�ѩn���u�U�JG����h{FDhNd�@\��1��/%�����X#�a򣉿7��-�T�JJc;���.�'a�pYzo@Y��(���Ҩ~�V�S���c���yq+�Wa�Rr� ���S���cq%�)�e�S��j�P��S
�x����1��Bv�V�ܰ���:_�%+}:�W��Ն]�"5�����7��ؕ�TH�(�;�cb!o��.��d��3Y��I|l����2jd���R��]�S�{���aD�w�)H=;�W�gC��7]1K5��u�|z5��:����f��m�7c�(�-�����t3�.���7ʻ���J��GA����40��x�>����J�#��:Mt��Y��V�����V<����<��w�O�;�b?٣�Y~͵���a�JH�/�YWN7_Bf5�u������N�{6N+���`��S߯�'��z�����7��SBGΧ
\�Zc_�A@�'Y՗h[V�7F>�kϦ�������"F��J��B�X˟�ɴ3K�u��X�u,�b=��;�%��HV��d��~� ����� 9�����B�{��:�E{�\�u��g���V���/o�%o����!�Z�͆c��p�3C�r#�5�����֕.���A��F�L�P�aB�傽�)��a�!��h����>_�]|��=�0��(_ڑ�����N�^�g[
� ��pc0}XwORʗ�Ҍj���#�ŭ�P�h�s����'�J(��7���%Jyn61�/a���>n>����{�V�����r�� <�ca�XU� ��okҲ-�*4�1��������G�c��6���HI�l��4I�3�WF;��9��j)ę5�Yrh�C�����-��T���<.�����O(rI��y$`�	_1`�T^�����_���0t�y7�����`�(�y�^���A����y(�"���0����J�Gp�J�`��D��C��F�
��?L$���P=�%�V����y���}�N�vѻt��n���*�;���]�C 5�7��ڣ��%��:'W�2�4���]͕B�Y�`�S�e�C�k8^�M���Ѭ�;~et�,�ڌ$�/Ň�I=��T�ľ�d��7a=�[��v�:��=��i�{�|p[��9B���ʟ[b��~�f�ji��`��S�tm��1\/f���<H�d��e��f}u� �uz�Fk�7*}��"o��Y�2�^[H�
W��<~�9���l�gO����7�0."B�;��<�[��:��6��dՠ�`���	 �T�_�@C�	۶�=�d��9�cA�I̺ ѫ� 
��Lʆ���f�l��lrT:��t$�9r.c�S��7&R�G����=����y5\BL�S����z[��J�� &����`�����!�Y�*�������>�PW�N{;�����i�=YA����3���e|���&�m#_�J�za�¨��t-�[��|u�ssGYLt�8p�%^����k���~o��:�K����.;w�T��a2=��*!���Q�V��K
��-�u�$`# ���?�\���*)[���?��p�^|�j~�Tb������2�����iϝ���������$;��eJ��ڈ�ة��A�<>�M7蝄��.4p� '4@!XO�l�ߛ+BL/t274(�#fU �Z_`�ot�$��O��bh<�ِ/�TĴ�g����ޝ��#�a�x�J-CE˱|����¹��tZ�~۔&���Zm
�W�����]��#�br��w���o�#6�X[oRJ�ǉc.�r��, n-�p�|�'};�k�_;V�(�(��tg�ƌ�N�F=�kf��3o*�!���ϣ�2�i���|�� -���k��.ܞ݋:��- ^�X��w�qRBe�)Lp�5q�YQ�nFc�`�̪�8�x/�YE������d�*�m��=�'�҆W���cщZ˔�7k�M�s�[�Y�	Hdj��%I�}=ɡ ��{W�dKp�q])��PqSO�HgYw�R�Yn�`�jk��k�S�d�܀/�N��_�Dz�q['�$��猾���}��`��h��f4�-z=i��b�E�e��Z�%�Ϥ���"?�����|��<��y�e��}�㉟�Z��gv�S�B���$.K��_��[/Y�j�$`��}A�Q2�'w5�sz�� D���ŀw��-�FD�ϻ�Z�����\���/�HM?�P¸.x�)�7�T�)��>_� ��V�I�;�h,PG@�w��]a��Mc��[�Ie�l��?fs�ÑrS.���2c�S�4��߀�.�ⱌ�Čm�G�qE2a��{�r��E:������x�%�O����v����>8o��Q�.�B��.A�Λ� �H�XM(LL��>	��Ɇ�x6obS8A��oݔ�ž<}B���)�i3gR���&�^�	g)�Gi�~(���
/��u�T*{�}h�I��yѧ񃴱�F�󻘾cI#.X�g�<C�n&�5���8�t��f�� ��v�r隤ة�W��7�"�l��FB���P��w������*�Ԟ����g��LB��J�6� h\��}��pR���dJz�I^�5��a�N
B<2��G�R�ɣ����yn�VN���Ѥ�rWA*���eX��h�8�����(�3�{�p"�,&!D4G���gce^�7���4=�[��	��t*/���W񦻂]�p�H�)\Y��Ë���~�/$���.�Ó��/t�^�1s���B�����Wփ� :�AX���"3�!�0���⺄����$>��%S�˷d�Ѳ�W�2U�����PK���o��Hk7y-{���4���ۉ��A�$|�Q0� &���Y.�+�^ '�O�	g�*�de�}!m��6�Y�%�9�w�Q��}���W�k�O]���K�M��7?��ډ �9d|px���fͷ/�<jV�Z��U��%}w%�P���D�T�T������
��$=m�p����k���m�AAFc�F��\np#���\+x]��1)i΁H�`��ݶ��q�-u��K徦O���R��27	]/�E��˻������/m���1_L��'��&��:�-��z5��_M���l�i��;T:���5���1:gD3"���F�|n>��Ф�E�P7Œ �������ɮ������p���RA@��3>a�o$H������l"��-�ӱ�F�}3��ݠ�R��ů�V��	��c7�$�7/��}�i
R}t�ZNT�Z�H��N�A����9�x@�:�f�����֘ǞJ�H�+_�e�abAP<r�4ʯ=}�+#������g������D䐊J�;HԗHA8�����L&�%�Ɏ��O�bQg�Jӄ���b��,�M�+#���� ��r����Ƅ�`k��o���:l�f[�&-E/�;m��8�|���P����>�����d������t#��D�s�����s �~C�#��N&���ⱳ�=��*]r�w��7O����l��b�ڒ��"�rp Z�	�<U�x�Y��r�|��b����[̩e,��g,�h�O�C�YLk\CG Y�pl��-����Q4f[��:Myܳo�l4(H�T��QY�)��tك��;�CD�:������;���ٵ~���4{2���u ��gM��H��OD@��U��#���V�	{��ޖdp��{L��l
9���&d�R�?��R���� ���6m|�E�[�296X7���9 r|�Y\p�����T��cMf���E ��\�#�;��nBhyz(O:�yu����W;e�Jw�7�9L���*,�Q=��~0n�9�=tG���=�
�@��U&�We�7
lD`%�&/�#?�P��'�Y�ʪ�}~����,;G�7���1��4��X�	+�4���8 �H�e��Mљa����8��`x���H���� ��g2�/Lí
��<�;1��|uc鋥B}tFG���W���I��R����M,�~$ʌ��э6`C�$违'<]"�O�Z�InrT|n"S��*B7Eb�"̐��б��Y3юX$�Q��k����~�v�-���E��ٙ,�]]�%����`C+p~�mO�����·�#�L,�Y6ŮY��~,���C�^�L��>��ai���&G�2'�З�2���X�/ʷz=���}F�M���F�8���E-����Hz�W1�"D�ѐ� ~�4����rE�ya� M	@�O�L��V*��$��DbK{|� �u���x�?3q��x�.d�'�����>W���8��R� Kd8���t���[xg�}u��L�~�⻑��?����jD�����S4�/�`XV��,����5ɘ�͛��bXP�-9S�Ia�DQ6��||���YW�Bզp�_���=a��L��jZ8�a������/��׻���<P�Ɉ�f"�Hv�,G�$����4�'�Q�x���pJ @^�Y���A��l�A7�Q�/X|ߕJf����u�),��"M��;�	�l�$6B>m�K���v���E��|�\*T�%�{��"&�Aj eٟY�1�Ξ������)W_:���1ww$ͯ���(0ju�#;�%�c�4ķ*wJ�Y�xv���H[����A��xx]P�U�3i�:H��Im�Ͻ��êe��˼>^s.�J�6hA�F�6�`�s�ܫ�	}Q������m�=�[���Բ�V���X�_�@A?��}^�s��A�0zm7LǺ]�^�!�1X��.��Qz�^�OF��/�?������;>�\�ΐ����_Rc�x��7��v6�`2���O���6��w����3��\�������6�e�Be<��ƂЕ�mr��w��e1�F!��"�E�f�E�8��-�4�,!I`K�$w	����h�8	�<9m<9Uu�h��-˗S���v7A�}qw�y:_�e����I�Z����Ju��\����+�\�I#�T�w}c��b��*ж� � ����m�}hwX��;h@ �л_���sxG��µ���R�����.��ܸ�����($B4�����![3�d�eF�"
@܂TXߏ9����p�N�?�tZW��n72��BU��#�����j��W���1Xb�r*>����4�wW��xT�aP�#ޗqG��w-h��ߊ��QҊ��P��Z�� W6����+fJ����`�'��ﭚ�8��w�"gp��ڑD� v���.�h�_��I����B[z��;e�T`s,�4��}�%m�{ӑ���m�(�f2Zbf
t�=h���-JG<�ʣ���L]5Y� m�%�d���PI�SUb]%�J-�qg�W7���)4QO!U�S�_��e2M&VK�iZɯ�WK�9��lUʥ�!�����6Z��`�%���ƺĤbD����@m1m�W	_C$�R膉��ր� I nrP|���~�M����*�LU�J"%�&�u_  4�r�V�8$ a��Ľ_���m4J� yd�{n��ND�N�?㺆��	i�W:�n��r��p�ZVi�1Z&��C\��ك���3�]�V�;�v7�񽗯���Ò���H|��VT���Bu������2u���W�fSB^z�Q�
���(�� �<Ͱ/c���2q��4q�j½@s�*(������v��C�T1�\ۅ(�1�i)��)4kB��}Ƴ�\�	F��R�9�j������X�8���@ѷb�����ѽa$�3�O���R�-�ӄ�I����%�y�	Ƹ��5�S��W���JW���ރ��2��q�eY��Q�0�1��֠3Q<�J2���&��mHϒ�v�Į�S|6d�a�:O�]m�B��[�^)�_�N���ÚL���+�`/�R��́*x�D5�h��s��m�j�e�\�v��d�4�Z�"���~�aI�Z��PCG56��J��,�g&??�;�+T���-�o�b�`s��f{�uHaD9kA�'xS�Q��Y��0q���X��x���)H�0!�S]Y�9���o|�;�Dm�S�T�-�Z����º�Q���9/�vg�ͪ	b1�^:��9z��pف��Nt+2��EZ+l�%'I"EE����L0�iovV�;f{�o�.tR�/|��$ꍢ:x=푤:5-���H!�GN�Wƣ�Y�I��}����B�mry�{1iGc=ϙ}�N��"	�W2(m��b�9Է����qK/nnz.�\w�S:̹0t�]��N%T��u�$y��Л���^�����"
�\�_�;�>���'
�&19Q�6�xH¸������k���Bu!��A���[�Tu^�]�����ĳOO����N���D�>.�؎��
�݌2㌝J�aY�7��}���S�i�iVtK��@C �3����Z�I��^���zD�AdYNUz9�mVn���!��lܒ��J��a�m�<�gs�Y�j��-�9%���X� �}�ΪU�D�N�"(�	v��]��FՍ7�N�Al?"3������ǯ̈́��T��)�k�!l��-�1�8���_D�j��&�<5�#�!=��Q�Cp��K#`����H&��IU��wFWi|>J�W���)�V���(&웡����g��'�C�j����#M�I�|�]�������Jz�����e����_U���^��۹d�r,�`�b_��mi�� Іa���Z�͝�~H�R�I;vi9��XCe��g$�0�.0R;[���HW�Ѵ�wV0��sH|Y\XH���`�Λ����᪙����x�KV����Ȭ#]$��n4��[LBعŰ�IL�J����;A���\�&@f
��5fe'�`-����A��%���d󶉐�brm&Ң�v���K���7h�Q ֿQ�Y"����D�g��Ѐ�����TlO���Z�e�_=ñ�u��@�9j�t��=H��{��A�s� ����w����`��P�I0
���R��1.t*�6,�V�8W���M��i�:	tNy���.���x\��7i|��3���Q�&���<�w��:�Dd�`���:j�@,�q����^�t��S�-l��X3��`t��}���_[�<<~�2}y�j�������+�����_ω�x�"�óӓ���>���Z�1�t_�$�]��9B%T7|r���]��T����%hd	JjV���Ļ��&��b)U[O�ƞ8U��bD�ϒ�+�b��z�U��ǐQ=��,�_�z��F\d��rS��AM�1DK�H;��`�#�Ci�"����i�ܛ���/V�o�� ?�o��U��#��=�'8�k�b�<�!��.��D�� ��@��B�5Q2�;n�Ԡ �y�s&�jwWh����C9����cf�m�"��k��$���F,�~d��k�S-|��8�'� @'܂r����ix;��HxE/Q������	3Ԟ�R`����I�T���d�ǃɃ��Ƣh�i���7���+��IT���S������� S_fv�
|S٪���'�͢2��a��t�����8��o��L4��+�߾t����~O����ZV�6ޅ�9����@��;.���X�tc�����Z%Le�E"�kQ���PJ�G��q�����/Jl`�U���>�n�+��uQr9@x/؟�������8�(����1 �!�I� �U���7-U&pq��]U�6�S�8Q܏ŗ�M0��<��{35ف�������9��Z��������z��[��3R�գf�+��QD%�0֕����<�ə���Ȍc'K/�h�|+�̲a,�<�$�>�H.;J�w��X/e���J����x7-0���ig9{ULx%Mm�(i!�V������أ�+fA�:����&�G�k���̑*�����긕�$��8���$F�
ध��U`mt`x�9�[�9Ĕ��uo;|u����r��7��{�f�E��S2Fҩϋ{�,���s����1�O�}��6�s}Er�49H�Z�u�U�׆����7�%�� �AOf�ch��)L8�cy$���� J5�nA��=�$���1��t
O���[f�aƙ�������K*���������6V�k�\\���Ҟg޵��`UՎ��M�M*ѲMQ$>��`�	m7�&�'X���əc�r�hǎ_�7���uA���?���Gf��L#LOD�a�뛘J��^	�3�BȊ�ʈ�ϻ�E���3�K��g�v6$7�AE��M��ĕ��Z�Ӈݫ�m�|�3��4�W�~n�Ql+������1�Lї~u���rĿ���u����"@�3vt�f$$����7�^=Ԕ)lbܮ3wW?SZ:jv�ݟ�,yAVr8�!I�����u�~�hl 0�Zҩ�KF���Zܵ�����/���و�9(�Y�0x�9}���݀ �\���du;;n����2)������%�#����J���8x���W@��fC2o2?�3�ݕ�������"e\GA=G���ӫvJ� �#���������gP3�G'���(��c����4`$�;ވh�����՟����8�%��()r@�e[��ӹ�3�?���R�.�,�eeu�4�ka��]�-� �T۵S�F��1��7�]�8��޲U�\�C^��)�6ļ�E����U�m�|�`,��]\��ϗU�Z��������b{*3��\]x�4�E��SU����򦒝I.ބ|xi�D5�
E�����|>ђ��r�.���Sr�L��o�.�*}��&+�S�g?�J��0)��K��?�a1e�K��w����j�3{MΞ�R�G�:�=�+4"���s{�cL7"��9�[�Њt�xb��~x^�b���1�����q���n[͛o <�I�^ć��@�����r)|M'lC�J�'�ڎ!Ţ���}�<�.oX�el��]��P#.{��(^�e�^~��Wː�b�֔��Ȭ�j�CK�%{�8@r�H�2�2����6)[ЗmLV�X�V璣�m�_��*�{�E�'�/ٹ�T��7��H60��/x$<�p�'�VC�-yL���Y��-/�̚���ov<�!v��1��lUu��W7+�f�Z(ޡ��e�����2=S������T�q�2;՗~�0~k��i0Y��c��JUͻ�@���Ǹ�U�nr�G+%_�jqK�H_�]��2q	��z#߅ޥ���Y(����NR�s��N+s�E/XM��Dn�q�����e&��ҕ���$��F+0��fy�r�W���h���߻���X�S9�uRlqƅr�>�oh���y��zo⹓�>�=<���{�/�z�pPNT���������y�a���:�]��多��7� �Z9�36/|)e%=j-����2��p}�;Y��#E�K�t��?���OF��ȅC����&����8���������t�E:���m�!��Ĳ�S���%`k���\�(���5����׉�Y�g��>@Qz�<+C���a��+�]u�BR���@�4����\�fz�YG��dr��ֱ�:d+�LR����S)b�F7�y�Og��(agU�т��Zt����&�gθ�\!���~7 �r_^��t4͡并�^��&������Hm5<S�%��)������U%�	��F��i���$S��"zS%�d���6�87`f�RT �E�jLA�����rˡ2}wZ�+�h��Z������c�	����ȧ��ɝ%f�o���ُuP'����U-�Hk�C1'{晄�X�4�g�z�9��qnhR9�O��?������7�l�\�gD��{����*�q �g�~���s�V�N��Y�DP�}��i�[��t2�F�R�[VS�c�L<��j׫�A��m��a7x�rO���(�T$j�E���J%(���@���@�_�y�f���t�Ax�0u�;cͶ��Mw_)�_i7P���e]1�ULb�&a�����u]��C��u���j~t;�Bd(1��۴�T�׸Dԫ^��jK֥\������ɨ�N��W�~�=+���5���8������>��i����pY:tR�p�0@�Q3����κ��C�	�y���`IǢ!	����%�~��v�H�?���#�5>I�r�l�ج�x�ۖvhC���P�����XN'���C���a�?�Orz9E���|&�-�]�.@��"�]f����/�6o2��]�B�
e��EB����N(�@��I����g���BM&�qn^�K$��L.(Xq�	)� ^����������/ܣ_镯��0�6��׫�V�^;���A�����/
Z/��i���
�1>h%��Kp���'H�J�pxp�M1���C7��E�^��4�L2�0���@�>Vd.�C�a3m����d4���8-�M>y����M}�6p�+Y�#���ܲ�:�kN�|Sҗ,���k��1OE��i��iK5�����>%*u�8���@�8܀���]�7�i�g�]OW�����_����e �I�GL¿��I�e����X`�v�ý�Rz�e�E�,C�?G��#���,��L*3or�L�o`�@s95G�sr!��|�%�A��g�d��_[J�>�W/��Ó6q�hi�Y�W4}��[��m�sю�>v#�<S+�dQm�gXC�v�u��ҙӀ�S�>E�5��X��|ڦ��O���G������L�L�@ 	�i�8 wO��lyDz��# �3E>���������f�
�
ʈ���� ��.b.ැ0�`ms���I�ǁ�ǿ\t��
�dv�'1�F3��������*���#C�U	O��׮S����<\c�#D1�@�d�K�	\�%�}I��V�V����)i9���j�ˋړ0/�~�yJ�m'פ�����o<��Ft
(;b3VA��m�JvO�m֗�ðl_R T��g�<?��S��V��j�f��l�3W�/�&0�^���o�ľc�*1�F-�4TP٭������X�+U�~9����ȱ��₶L�#�>�Q�K9�� �\/IF��^��Ҥ����&3���w*@��$8����Y���H^	ү�t ����0$ǧ,|�p�FGI�dg���"�oKG���'X!���&x��7F/^� E�J	��蒂���#=��ʪ���ud0,�������v��Hb�o��T��hIt5Q'�YD',F�6V~ʟ�B�-����⑇QT|��@wS���ww�J�<�½Ǘ��#�@����R�	�X@����L(06�R)E�����^�j�N���>�F?M��m�����#E��0��)ND\-�̙�K��.�g4}���R%�����Wu�w 5����>����R���7?�R�")`�/e-��ǝh�d��K�N� Pr�e}ѫ�39� �~�6��Q�Ȝ1n���;�5ߎ7�M.2��(�����h´%Ь��I�m�����|K�W��Rt�?I��eYn���Ӳ:z��,'=	o�T��9�F����?�"�.9l�]�t�w���=lA�[E�r?���=���/ʡ����"���a	Z3����de^�W.�� ��R��p�xF��39=3��S:�'c�h�̶ݻ���{��Gn�oT�ٔ9��+<��u�]��̂:A[��|7R�U�a�I���]�jaЖ�g�;c������{�u�^���u&Ǆ�5|m�����l�&���/hgS��4�������F�&"b.d:����=�[oX��ժ�����~x:�* �b��W�����@Q%�엪L������vz�+�u��}t�����4�g��	��bһ��\�&7'N:�n3�C|��dڮtG\���a:�[0��y�H�χ5�6ֈ�h�-<k��_o�m�7E��	���
,&M�n�����e�S$�� �׬x(�-�R����s�YH}��_�^~w#�Q�Ag!�_�[ӷ�����g��wh;t ��0����I�^O�^�lM=\m:"s~���R��ۘ��3^<`xl)B"��;��a�-�R��W�8]��z�p��8���A�l9lw<QM�H$F���Qrq��U�� v��D 1���K���1�c~m���i�ە��O+��k����5"��'�A��J%hA
�0���WRXR��NA0��f�X�VËF�B�l�F��g	n�������FR}A�E_˄��Tѝ,�i�p��BZ1��]��x��*��yN՝�ɽ��W�0�����K�=XAw�#j�p8���}v�����gKH=�PO�s��hgbx�Ork��\�uQiťR��� a<��߾"�����j�a�˝����� v������i���X��e�L|�T��r:,����_��sn�D�`��%���ΪG���{���P������+�rP�5'� ���j��~�}��m�S���}嗥��Z$�7��,�PE�hՒ��������N���:���H�|;U`[Ȥ�ך 	��桮�5M��9��?�A#] �^Z�=�P���O7%�@
�j����,x�{�KZg�=ڋ���OGzy밓i�t������ul�2�g��;�����x�?~�θ��c�:ˬ�8t܂�m����h]�	�\��/2{�z�S5pr��weU4��s�"��o��]� �i�k4(�
�F&�d88M7�W�/i�4
��ϟ�VN8�f���
�7i�})/�W���TAg_���_��+����nT�qI�� ���MH���Ux�(�������K��5��w ���(��~j�f"+�xEE��u�
��mQ6��g'�	1�ߏ��H��*�[}��QY�ۭ;�^��A��';��
~�h�LHk�Qxդ���	��(i&��:,�S?e\U��A�F�M{Mt�o,�dbB^�O�*R�t	2��:[HMxձ��L��
]D�Pݐ����(_2F�~$Y ��+*l�����ۇ:\��]��D�~u���9x ��&Z1�;-�%C���x?�1U4F�j���M�l�:�Z�T07����}$0�ٿ�Vο��x�%��M|b
��@���{$0�������a�A��πޫ~�&i�.d�V^,����^f��)�����"�'�L���ek��U�`�4�PB%�	uם�E�6�p^%�Y�D o�~>a���٥�2=���4Z�e�HG�*��B�lNZ�7k3).i���01��7�*-���[���ӻ���׿)^Aَ��v��y�?l�F2�a1:2C�)���s����)�1Z;[��+��!�.Fe��}>N�C�ד�%�Ȱ� C�V�f���y����_�x�o.���FN�!�lI}_Û�a��C����~�{�[1r�0կ-��B�5I�N_ؐ����G�	�"?g��ٙr��j��d���K��T��C��l���XU�n@y���3��c�E�}��>��x8��u/����%ҋ��XG1��_�`��s_�?��i7�Oz	T?�^b
����%��3�����$�+���匲ŅW�ꨒ!^�C����"��"�j0B�'@�� �eUN��a[,�8'쨈lUM��`��E�P��2i�ε.�vcۼ���+���D�A�;�k������ݨb$��n����T�_��%�+�b�f_^�/�f����d<u�Ռ��8{����w�sz�:Y�����7����������eq>jn]��l���;�l	�g����*�a�>�NL�4(�=b^�Y6�)��&��^��$�ì�	q�Kt7#󲝅X4P�/�T��n�|d��!��
i�G�"�3�p�=��B#���r���u���qY�:J��Y1 n����ː`��
�x˙v4����h�X��,s�w����]�g�2��ciW�Q?���"��d�su�k�$��z��qF 7	�8�/�]%�Y��f*��������?Z���w�U���cS����F�3Q��ٰ�-E^��1�c1e��H���q�Z����:�V\7�B�J�|���q;.�"#��0kC#�\iVU�!���HF�WLI`B���N�?K,�p[�!�^�j��w�KG	͝��[C�'<4���A�ju@��mdlw��6>֛;�k^�ܟݰ�	���<�$����\\�>�����P[�w��F��>sH:[� ��
�������~�� v�ND�?�j=R.�w+�ܩ���wi��%��KhIڹ���+.7��ww��K���n_G��m"�gB���B�vg��kW�uOs��ۉ�.@��!oM���� ���v��1q�W��Y'S^|L�G0I���h���C���.�� "���g���P�[�����ɺ��![�W�oX��6o�Y�C��T�0}�f'��	}�V����g�'������;RG/
h�/5,~��0J=�;�>I[��-�~�:;�6�@T!�!`FB"��_�6�D勰�*��Oo�U�=���%@#��p�mz�Ij�r��ۄ�a�<]f�pm�Uz'�`l�!�B�i�A%���BR�v�E��۫퉪���'��!�Y���,�%���BY!�] ��Y�}:�*�#�Ɣ<��.�?Z^�)��9Jz���1*�.�?����77�?��b>��?�m�]��N�c��HɁB�]Ҧ���^��X$M��W�[ˌ3ԛWD��AR1=�C�p�cَm>�%�/|�./��s�<#X�ў�����tX5�>�iP^�N�V��1��+��v �/�؝,Ѻo�dsi����4Z'�-��Πq�nAy���H�A�m�R�^Y`ۭ�,ad����@^Hv��~%�O�w�V)r�u(3y�[��8&�E-�B�'��-]9I��0�XEp��w�]Z��-4t��(�D�(//x��UӨ��XOP��~"l�I��Q�T��P�X�x��{_.��l�K���Wƀ]���Oۻ[g]X&�C�]����އ#+�_["��i��ǈJ�7�DIg4˧�&�%t@c��0�[=�����w?���Iǆ��b7ɭ�	�Gʱ��'�1�cO����s�tK}���!�rM*�aPT�Se��[{��`#�iz�͵*���Ryi���M�"唧��e#)k:�$z����4$ݛ����t�AAU2���Gǣ>���z�߾_�<��l��C���x��٢�Q=�}�N�w�$F�&��\�~�.n�2��%��ߧZc����#��d�7��@�{-)�Ќ-N�~<�/Q�	�"Gu�����r���7W:�Z-�[�����hp���C3�����qY��&��.��&>Jf'��k�d��I���&9�m�--�kjU_X�2�O(�?+�T��"ƴP��.�a>�����v\��1�o��w�웗�~�Ԅ���7s�I�g���u}���+�F���6 fxP����VuD�3���DVt\"����Bk(*�~����L�X��?$����̑m�������TW��vh��i�}��i�c��l���~��:��#�>�vԱ2u���eK��9���3�І�J\���l�9�o\�l~�C����X��qn[��M���s�vQx���qp�1�QT��)��^��gI���n���X7�݅���΄~ƴ�f� ��k�͇#Ky�����%H��J^��̊�<����hR�]������442%��ԌК����V{�
�v����8�O�?6ty�L�R-�A@+E���y�W��\���tܭ��U[-����]!?M ,	eϓ_�ђ?QH�<?!�}���.	�,H�MV��m��2���-H�\�a��d��`[�Q����F�����[����-.�0���&�o���v�nsm�H�?��>~�5CJ�> f0�s�[����k�mZ�U��c��%�����k�������nk�%��/VW!��O���f��C-��3��
�zY���x&t{�Ƃ���������_�Yh"����1vfޯ܈��`Lb�c�L�kٲ��B��J��	���/=�������痞��_cb��������WL�>��3�!h��Z���I�CX�}���'jid�@LwFeM�+� _�xN)^�ͩg���	y^�C�V)�j���k������g�����5b<�w�|`�|�a�ۤ�r�N��٭���1�ь���o�kA�j=1���
�u'6""i?��#j�B�0)O���W� ����( �#a�{(��Mx�֫�E��`�b��I���pf} �I/�J�Т��4e-�w�.Q0Ak��I+�Dt�HWvP:�l�[�,-(�nD3�L����1��@ k"��g�d�7%>�e�r��q��"����D@s+Vd��d@g��Zk_��C� ��|����8��T�Q���c���g�n��y��x�M��Þ�0�l��y�Xv�s�,�D>��pG]�$����lٻ���ʚ/��w!mJ>�R��n����E���Q8�[��=�N���|}��yl<����AV�s����@�sjĨ|��n;�)�����`��A���^[W1N禧
R{��:-�=�c���Q����Y��O��7׼�؞(V�a���h?eY�r�����c��s7bL�k/i���+��3 �vSm����6��PBcr�0%E�ߧ<���6[���������7�6�$/�<吠��\B��3X/?k5ư3�ou��j�%1.�|�)4���=o�.,h�<W!$�#��Ū}��џ��$��C�#`�&z���%���P\�U��� ���f����\��}���&����9d~�ƽܻ.�Y����я�QH�����F����,{�a,�m	I�sl��_���RN�>vV%Oǵ&#W�\>~��Ā������l����؞q�b��iw;s,�¶�i��7���>���h	�:D�4����G�$�AZ�+���]�*`=��d��񸮀gU���ԣYurm��R�j�US&J_�-�����&��m�|���g(�D�\B�g#?�5����ՍAk��vt5v���mo
�TƓ?< �A�.��R��z�䇄$Ym��!D2㈉�Dx�]V���E͈V�%=;Ih����I^lɪw&�!��J�n��?l�#eo'M��p8� "��2��&)�j̳���]��a<z0<h��W��~|B���8����v�P9~�`VI����i=�)?�-��ݕ��28gC����d��=�Y�z�mw�8���Sc� �0��m%ղ��vI��4��+� �؏��{y�e˖q���*�KyZ����ޕ��ʝ��mH<���8��]�h)P6Qڬ@��r�3�a����6����1����.��Mc���Om��
��Һ�
��t��/)H͖�M�EG=G��j�L]Y/lF�K?^���찪�t˰!-v�kt�u��kԮ.t&�▇9S�Q k`�~P����1 RYN���J�N��:�I��t�"��m��,J܎�M�̳|��j��[�w%%~��k�v��1Y���'��Ok/��ǯ�#OE�y�mK`u/�%�mo�"�k7��!GK��P�؈!�����Jjj%F7�3'Sa�5ī&��4mE"]f�X��|A����␟��Z�w�c�d���]ua�4붚^g�e&��6�0�������
\z,>e��{r�@A���p{�;�	�;�o�����]
��j��O�r9�H��3.�~�^�R�;$��s(���!�횞+j�M>n�� H!&�&�f������_���8�-:-L?� iP_.�"�<i�=}����[U[)�ĘC���S��*5�{Vo��=W8�4�83XE��g~����!�|����r���k�@�Y��qW������?�,v�y��]�?Ȳ���@-��$�����_oJ�U#�7:;Kt�>���B�@r'&G�GM�z���wn���>Pŉ:�o�n~�	���� -�z��g�m��<����:�i]��bN4��!xZg�$ND�`�n������g�)�By���~D�0����i�
�?C�lOB�>x`���G9�ki�~8�hY.j3�1�SE2s��&Ezx-�1�L��D}� L�[6
e_��|B�G�t�A�WM3z�;�>�D�[��M�$�1�[�mȫ��Y�~;�g����X^%t�W:8(����9N 5MV'e�}����qG�Y������&/�r���m?/��1���۠�xS�d L��\�ɥ� ��j{��1�jty�e�Adl���W$in݅�V]Gm��l\�w�Ćd��~)�:Q�H}V�AxBV��w�~���&��L��횴�!d�r!�tn��3�թ�bb��H��ot]��X����t�A���_�Fr����!����-��P�Cj�*x�>���崏��֤k1�eJ���8�r�%��-��C'|���ME<,Ƶ-�I�=�/��<�o&�~�<�q�)IL��6��j��������T��]<a�ƿ�X�	�ej[�@�2�G�8"�f�O��4�G�Qz	�/f&�,�j���f47ܵ6�j��ÏWpF�P��-��{��{8��JG�t�<�� ��t}�Ep���\�g�3s�ɊL�tt�h
g����77�K`��C��l�K�٘w�s��k�o���d�	$������CJ�uuX�d��0Ó���J79�����ډ a�h��I�p[d���l�6��g^���4:x��]Z4����nh�i���0l>��sS�*�<�B��[��7#KNPϞ@r�ޗz��G�P�Q��4'��H�I/p�`�9/"	`��RE�&�g ��K� v�
	&.EM|��q��?��:�ˈ�I\��V� �d��sҩƧ���(�����
�i����0P�����0�}�ڞq�O�J�l �
^�P˩�^Hk�iv��+x�AAo�u�7�b��t��c���~w�T����aye����z�W|�O�:e�3m[m֨���J(��v� ����/����͖��0K9�Agg�z
���%Ɠ��ސ���"i��M�j���OOAka����!�|���n �4D5t�Lo]�'�a������dT}U����S ��x�(x��W������ʡOx +C��C�S�%��������b�od{ŏ�+�q��5���*�'�3z�?hҝ)�XSA!���t�J�aFpX�3��g��dQ�~`�e��x���mv��������Խ������{�fp~O�x)���s,�uB��Av���E�7jZ�,Ƕ�;>V�bԻ��'b�5���r���
�2F���0��|3������Z��MJ(1k���'1(us�/VY�=��[��%�];�h����5*��x>�-U���k�n��u����(E
��-M!�=��i"���bpr��L��
�q�oRn���9)�ވ�7G�ɒ�*�}ߣ�^]��ed@o��m����3\(��\��mK˼g�}(�6txQ ��j)�׽������g�P^L������g#+6,�=���G���懁��c�Ƚ,�Ia}脀N߇Ry��PG���`�����u������Of�}�{�.f."ʸ�@�����AוH/R/��5h�A�{rB������<�8��ģ�œ�<_^��'O\��
[��~�1\Tn(�C����/H��g���]����jE&gN��/�[�B��i�"tו磴�M�s���_k���u7�S8�]2�~��d�%¾=ȿN��<��X����
A�lY��Q/��S������8h��Jj�S��:��aF1.�چ��_��h?X��"�j	Φ����ͦ��
;�x�>T��6��rw���M����a_���	*O��R"�;$�
5�s�-y�h�8ςo��9�v@�i��ٳ�.��/�Z1�t�Yt�_��CߌlBU@:8޹�R����Y�0��^�2v�S)	�0�f�=M�%���НS�T�V�\�t��o�:����MT\!�C�BU��y��'^ܔ��������Z���v��1��h6�<(-��=��[\f/�#Ϗ1Q�§��X� ��ZnW|,��6H��4��I���a1�Y���m��j�R����>=J��q�@��_��/���w.�(=���	�:�����")LLWBOJ�Hn��AT$��{_�����D�;-m��=`�둃�z�������j&�J�g�g�`cH�(c��E�K9�{��z)p̬f?τ�yir�� k��$���CH?����Y�����pU��Z�=K�<����n,�<�=�3>�U�B�3"_7���x!	���V��"ܰ�������p!&�l�1���/+v��z`O��Pbg�"4�}��ѭ�_Ist�T�5M'�n��^�E��װ����:d&I?)���2�(釷�F��\�U�sk��o�o���y��0݈�a>���Xl-8��I�/G�̍�H�f�!��k���S鋞*7�gK-����I�nn��a+����:��L_���B<�do��i.��p�&��IINe�x�r�W3D2dc���5`�3Lm4*��r�� ���)���I�5*j���~��7G$�01-������ʋ�@>Ź =�%v�� �%���b[Ð�+���u�������O�r(�5�!���zV�]X[�;�ʱy���o�����B	/,o�-��ix��pȡ#E�*s�ͱ�c��R��\z͂�T�� M�"�����g��V��e�ᝅ�b� &�1����R,؜u�Nv�2/������9-��?YO��Q�?�V*��x�����f�Q���J$���Wk�mZ��阘G\�4;��^�L�6���Z�8����2Nγ�A6��z��3H���PE�ؗ�-�r��{���QQ�([2(u.��x3ޜ�n���|b1@�����uϘ9���[�DՎ��E�4��:��\��<g$�p!ev�&���hd?ƃT�<�D*��(vJD<��D*����`��������oSl.�p3�j���>��DP:R+��$�-$f��N@�9`Z8nK5��݆8&.�x!��\B��XX��(������Uo��>8�|�7�A滶�|j}����
.��K�[G�e��j���T�9{��J�"r
�}Pn���,�eV4���h��e�9�65��T��J"��y�N�5�����Ȩ{�P5{c딧�-�8�x��\W�ʵ����x�O�>&��rk�
E��]�5_j3D�������Gci_�r'�~��� �8?�z�r4�zꀧz����R���f	��֧hջ���wa�� �I��OcW���1>�q�fdSz���V�t�2�!�M����?����]oE�i\328e�ț��^�y�T�yB�]`uذ��w�d�>��I�{~��6�bj[ۍq��[s��{�`5]��T���<��
�嘕:١�l3d>�ty����� ��<4,������>QE0��9I~y�#�v����6���c���Z����;�I{�Y��ղ�����Юq�|b�Qk�BhF�f�,u�g���v���L(�5 (R�%�s-��^���@��[�����^�������Ŧ�G�O:y���r� ���j7��yT���AwXMtH��A�wD��j+�c~�kW�/-�h ��1A�ׇ&���t�
0ٿ>��v�%)%S���.S%�h'��jM��O7�-�~<P2���:�YƆ:�)����Ëe�"�ul 2�>:A�hN#M̸��?��'�Fy���y(�B����td�����J�BՋو��S�-�T3���[�
0��U��s^�V�><2�"�4�����Ic���E{4�Cc?��.Y���ߪks���ސ�Q����X~!wWҀ{Q�9H�om�[z��ţ,ܟ2������H)�%=���QO\���q�y�Ҙ)גm���fj����jv�\I����GB�"`��jB3Nյag4�n�h��.��nF��:���1N�c�. )_!!($<$bm1)�BPc�J��˓>vx1�4�F�D����)0�F��n��XliO*����y��y�!�e�9u��!b8z������ò�vËS>s��W/ ;+s�k'�>J���
=���"�~l�h�CQ�G������f���2TJ��/9=�'���O�x�o�JOwr��<���o)�zK���m�"#�'r�Nl:d�2M+�8G�MT�^��c��(��+����@��'���P�{8����Z�q�*�5� f���{�tN���~���Ȝm_�� ��#�Q @@HqJ��@�.��V��w�*oՉk�U+����M���FZ�h�]�I¸lX�޺��D���G�^��Z��|�_$��#��_u��������@��!-����He{��$��L���d��������	׹��WԺ	KܠMU���χ�ʦ�C�3�࠵����maZ��<"[Ʊ`�oCX�Iˏw��5ǍC�t㦌f�j�,K"���Rx��P�HWS�ųrU\�+�{�����=}"�[b�f4�t(>}�Iz��*)��+�,��x�2ț�ǋ���NFK��K]�z�Ǘ~&6[׻�ٜ#W�s� �c���_{uS��EkهP�Q�0'	[pR��e�E��׫�+0���6T���H�K��� ��jG"�Z[��u�x��!���w;�x�������Q��|�8)q���ѫ�K���j��r2a'y�Yѿ����V�a&J���K�|o���G�t`�\���IRs)W��PpE	�U���q����⢿��EZ��	�{� ��xՍ(���m��E�T#z$�o�'7��>C���������0�(6�Q�V�r�r�H~��NG�o�E׀rRK���Za����w8
W���)��O-��kO��\`Љ��.�)��.�-Q'r[{8�#* �-	ζ��)6�W���,eE��I�^k�Q�;��EC�p�Ѻ�/h�Z��x8��[�#Z�Y@v0��Ð�Lae�qu���.�k4�_��$������36�*�U��!܅���	��Of�e�� ~�.e��u�+�D^�]��R��Gf����M!���äFj���8-�V}��+�w��j��j?ٷ��ܺ�tϋ�P�C�Dѕl��c�ۏ�+��R�Z�T�^Hw��L�������R��n�ejM������T6���[� 4쩨����B�K� �R[�m?�C+��
��i�1&���kk��s1C���?F��� �ߐ_�Zͮ���u޼HQ)e��ـ��*>��l�b�x؛Lnҭ�ZD	�s?H�h��ZQP���z�����-�5��*�neB��OB:�|2Qb��/���O���h�^-�ѿ?�V�9��������Ƴ�"q!���Y����hF2��,��"��Y�`4\so�	�y�@�o��]))�S�����pS�먏�g�ζ��O��P��h��h�(��������E}���*�*�����{6�bÑ�P=.�^��x��E͊�GL�&bM�A\�E� �c�T�?��N�"��eD}��`��\8�L}#o�5�/Ӧ��+��\I
�=��RŻШ8��ȧ�z������{~��kwP$`�p�A���K�X��D�o��k>N;���O��\��{{܍o�����Z��
[���m^)1��#�y* ��X���j k�}Q^y����C�`�Ϡ$'�HJL�L ���0~5��D��C���i�Co���g�
{)Jt ��x�P&�:�Cs��n�w��U��� �E�$�������E�����2�K-K�>���Ԥ��f�R54JT�L��l�~&5Y~��A���Ĭ{��D|w�Q�1������T���O��F�6z�3�gS
��
#Z�d��P���y��6k���/�Vq^�G��wo���]@�b�gM�O���!�fnsU�.,x�]T��B��	ڼ��B �:G�X�]K��$2�X��O�^`�B��7��v#�V�ؚS,���Ձ�2�AOG����\�|y�DB��r����O���y�6�)AS��2s�) 'fƩ �M�19�Р�m�VϙP��Ff�4�l;�AŢZ��;h��<�}62gn�9Ɓ�v�D롫��kg�X�nA3��ߙ����~�x��������M纔�^�8�>P~
�	ճx�V�5����`�[����	�J��:���P�'r�j\axX�s�J�)��*uA��٤����������`Z?��U̡�K��հ��V��+U�v���]��u�=�B�K���F�4�
�_�Z�ȝ��>u��0�~��|T�����l�m�����#F��`���x; �S@��`��q�y�d�4�\���C��#���rꊫ�^��x�C�s���y�F����t*[O$̛�@�xv��?t�z=�������OY��s��n�����B>R3��v�m�,t��oY�3������|�������<b��/�19�(3O��!0��P.2���p�n�v�[��� F������J�����ݔ�I�u�q�A�d�&`�<�U�s=�?l��
\I/� ����Z_��b)/TM���i�h���fJ���bXg���9�+��?8�/.�A[�[~��=�}��ж�������2Z%�'���P���l��5 >��(�<@�/������-��m�s ˁ��υS��$�IF~��7�������!�X1�x��e�=e|�D�;޵�����+�ws���b@��Mkjf�s⾍W[���cҫQc�*�<�=��:��Z�x�\T��V���&�*"�l��Ȍ��v�R�U��i�ֽ?�*?{��ð���pG0o��i%5�{��9t��<���[-�g�H�_K�UDSN���Ԃ�A��Q�{�I7�A��K�y��T��q@�e9�4J�4�q���z0MM�@#m�c��;�\����B��E����g�r�1�er{�HlII,~����N﵈[ŁBZ�V2Os�2�sU#;�A�n��[��W���,�ޓ,�V�������Q�[�tŕ�Z<�ø܉ͱ�T)�>c����}A[�ޡ�i4��~pm�aQ���L�w���bt������'9����Z� �&##Lrj3�Хc�Ƒ��V��G�,�{u�_�:�� wGJ\�.'�m��\�¤\OqJ�@����a�~㈈� Z
��Sr�v��a�8�U��w���0F[l����>�����L��+������⁣&���;s���~X3�ו���ӯx&Wr���r�/S��z�ҋ��ֹ�&LkHH�Mv��#�v��l_�Cq�HO�!�B!5uD0�d�
��\�8�F�(
;�8����QAJ����ܰ*���t����#J��M��7AڱY0~����MdJ#G����r���O��y���2�c���G뤷�;5.Xj@x,&B��~��}L��ի<9��?�_���--ٷ��F?g�ay�h�fz�];����M��tY���&z���v��Ѐ�P���6�?����@��gr����ZQ�w:�/y==��jD��Z��Qm=�x-�#Tw\:�~��� 9��@�JR�s����)*�V�ϖ}�e���W0�J<��f��R|�3����J�9�=��r�(4M2��\�ڌ���)��eV�)���:Ǵ�;�Ңw��LB��:����,4R��q�v1�s�Ͱ2/�J�������X;�Xp���11	@�	 �C�0���9+)&<�n��+'߮�����`�i�/�۠R-�k����Q���tA�(�����Ă}%+e�ޥ�{)o��q��J��E��=�c���-�!�l�B�^:P��3�M<�j%-�\61;�%��a�����H;x3�^"��T��|��Ϸ��NQ��������ޘ�.�Qg�&��v^��,�2���_�F�~y=��[��G&����B�ӷ:�]O8'U���}����؛�֤��Q�pͪ����W?�3����/��}�i�wF�����W&OG��DAk���ڄ��$�2�E_�F4T^��y~�����f8Ug�|�7�!�xY;X�"oT#�{h��$@�yx�ꠝ��v�:$h�B��^���z[O�3=�Š;��Q�&�)���������o4L"������v���[�t��� \�{uwx�g.hA�%��p"9�>]c�@��
��h1)���/�$��_n/r�ω�!%;����ֺg%ı(+)5�f*/��'��X�I虦���aS�T����e�ɒké�^YH���7��Yg/S�~��^O����^� Kh����,*�޼�L%����X��vjT[�ꦒ��罤f�F���F"a�|"_�:	?"�_Dlzf�i�r7������u$�N>���a�wf�J5)���X��b��TX �m:�&���13�'D47U+�}��i��5V6�$�^� r&]b�X���#c���v�1�*L��HH%����7���ḝ��~MD>�ҙ���ߜ[Y[�-	A�<�����!�����z�F�RBL�>:��3y�Xj
�[���e��L1�%���F~O<��~��'?i�����&Lx���cnN�����'$S��"��w��A��j�g Bߧ�t�F	�cXcE�'�jS�s��R�.�����?ܟPMϸ�eۿ�g�?\Jb�	1�a;T䐒��b���q
����
j�m)����J�-���w�o�n.��N��-k��x�"�����M�9a�z|�xd��;d�h���laω ^,���7����6� �*��������/����)�`e� �y�eY���%l̬��;�u��R�U��+��$���?���CX�<#�A�bU��X���H������l��������I� �sT1�^�^������/��X�l��D"�)�1-����dG;,�Pe��b��NP�j���Y�ۋ#�b�Ư�VV���?j>U���ͫ�9Ie-���[׿��7���h����RC��������E����Ѣ=�e�4u�8>{J�,�Iӭ�r��-S���͙͂ļ����S[����h�S<��Cs�0{�xgWs�Nq҆,y듹s��!aG�::L��������w��a�攋�z�8=告��J���r6sD��}og��s�V:Urδ���h	HM 2KA &��U���/��W�����gj�@���@�mg<���c�\1F�&�lL��'9�$?�3i��q_�"�3�֧�ܳ�x�U�/�:hKV���ra��7�h���B)M�b5Ѐ��-j��]�ӗ�'��E*���E�zO_�".�1���w.4�K���W�4N���a�;�Sz_v���Q�h�E
���K�7[�q;�<��������߿�	�������Ʃ��-%��/�g�J(�����yi�p�m\����*	���|�h�mˎO�^_�Fa�Y���ejW���&LO�p�*B��w,��e�D�P�Î�!,+����j��t�z^W�489�����2��e Z{��'�.ə.�xC��	HA��y[I`�g`�c��'7�M���F?\�/a�i���FG@�D(U5�P �����k6)2O�f=e���)�a+�B:����J���q���.=��/i�n��K'�]_9��CM�Omɋ�@�p����;�Y�P�tB���ES�[!�X�h&+�N,M�a�-�%+��e������u�Rx���c���|n�6�H=��v��f��)��3 ���5a�Cl� �HNhB$�+��B`u���9��e݃��i�,�ZK �����"�������{�c��IT+��)H�4����X�v��9��Q)@j�z��|�E3u���B���Vd�Q�G�:g=�t�*�(�R����M�	�(S����Sܫt��9�D⮨;`Їr2T�H� .��7R�2��Z�z�+�{�-}��;�l�t6�k�<r��F��'qw��VT@R!���5c'�k%��-��~Do_G&��6���NѺ�}Rr�,10��45K��J����VT���!�������g�6���D�~Z�#���+�/�W�%n��ZsD�7�~ �{�,V�YLί�+n���b��?P$}9V{pO����J��#T'�EoP��T��
���6cs؏�`$h����PN@S�9��C~��`ˑ-��Wa����.>�*�.g3#)ȗS���4R�ؚ.#*�.�[�ë�`Zm׾�	y��]�<��vat'OܧO��m�f��3����v�ؿ���q�}~tZO3)�6(&A[�M�JU��s�~c��1��nG�-Ur��}��ʭ��"C���P�eZ�!�'�ܩV�X����$�p�O���c� B�����:Gބ�q��i���H���'�KA�!7�Z��V�L�g�R��V���_R�|6����%)�g�Q�Μ$&>�+}m���>W���a��\]r{� )�\Q�v���>���Z��h��8���0��r�y���)�>.�4brs��*���]�r�ӭw��Q������|)�7E6��}��Y5;C�L��2�W!q+S��4N<������(j� �A�lC�A�us]���W���6đ�3n��.em.Hg�����5T��Di���\�(�B���{��_-1&4�����k�C8�������~֍��9�8�fv�� Ct�n0�X�>w@.X�`�k��0&��ύh3���:�0�e�$n��{b*X���n�)����h[G�q�������ӘI��c��CD''���EdR�g4ZS���>b��0*ఀy�؃G�������_�S��u��W�!���*�crr�0'vn��0��u�*�^��z���T0Ų7q�\Du�����$�3��@e�)��%�(+ۈo�e?v0�����eÑw�(�z�3��'����Ԉ }���Jh����|l S2Q�(l;��l�f]��=�k Z�Ʋ/*�$�]ﺦh����1��&N��}�?��������q�6� �õf�>R�k^%���_,	�eWu�0F�N*>}��'��(���:d3�*8�*9:����u]qc����kwUn����1�!�H��P��rvAA�ë�Y�Q%L<��?+�_�m�B3%Ye}&�Xی۴;�Ǹ7��*��ƳӵNPD��������ԭ��4l:չ�9b]1���r-p�l�Q����b+0?p���*LBpS�V����sI��r���%F�Z���T�Y<y�'?�����}��}���!I`���>-�/f��,ļ)�)�˜�jt�U���Sp���k.3�s����ȓ����=� ��mzD�M4r����c�=!���|���d+�maV����H��Ldɷ�F�8#%�@����֦)�.�6��v.yޒ�U^4�����=����[v�yё(�d,$��_���������%?A���9�^�F��sfߵ��0D��K��bV�^�C�A^�\��]�#�_v%��D*�`P�Z�U�KV�r����T���3�ß2��ҡ<���d�Z����Z�5I"��)-���5H�H���`f�c1�����*"z���z���3�1o��;�e�B^�4k4����O�&H��N9Ҷ(Zz��.� �uȃ��ؓmWC�Z�N��MZeL�� ���7�/+��m~8W���$M�ù
,�ʖ��-�?_/2]tJ�-j������d��5�n~
��`�*%��mp�'G# h�X�}`��20�Z�0zR�Z#\�>Sj#�G�i$۞�2HC�^X���DL{c����1�{/Dϛ2[���X�WS���a�W�DШq|��ީ��߯��Fl8�2$l���zp��OP޺%���X�p��d��n����!qGw$�W��g���s�7R�6�2�����f2N���8�g�mMv{��H#DO�1o���1@5�v��7	�~n#���u?�����b����QC��34T!�n��Zef5�+��骑gV`�����|$���(�֜	L��~o.��Ɉ��)_�!U�/���I��� bV[Ȇ�R����H�3�1��N���ؽ�6<�Hl$�
�|uD1�?��DH���|�1�݅TK��%o8���褓bM���L�v =d��U�ҒrG	MwD��
�Y#��=���,�Q�+���әR���'�R}����e5}��E��-�Z�T�S6��W�D�i6���n��z��l:t���xze�S�ij���"�8WY����a�v�qc��f3�㛆�͌�QR�8���8k^K������_W��K��=�����7g]��he�Hcσ����|^�*��as�k���뮵��U]�fb�,|��F.I*�\Y|�13V�Л!�o��s�Hb7�p��aʅ��R��і@	-sA��S�ŲV��$9�~M�wQ��z�g��}YZ�s|��&��$�$�槍x���H oM�4��?�!m	��6g�L�R4[g`8]AI� �|�Ю�0��f�F��%`I�k�=L�'�э�e��)��_Z�Y0� �	�ӹ�^��SU�ט!fh�# J
ui�b�����+����TiA��'��2�Vo�~�k�U)�i��,'��y����u��"�c=?D�����SA�I/�-��\�����H<#��98`����=<ȼ�I�yY��n#�����%�y��r=|R)��͌J���4�ģ\"�RU�J��hzO~�nA��Q'I������j��pp벼����}��N�S�Od����`����u�&@�83��� ���/��3Q+�[5�K5'R1��L�egፉMK�0q͒����Arw���� �W+��P�_����g�ssX�J.iy��"H3�jV�b`�p�&����v(x����Jۛ�H��ht-�ֲ)�f2Yq��U4ϞO��E�Z?dY��-/@� Q?r���R4f�y�%=8�(�qQ�T���sɣ_���c�� U�Sg� �F�f]ӣ���Z�m$���B�iE+�DV�]y���]���)ѕߛ5s3q�ɧ!�VU\0��.Y�t��#Ф+Աo�?������V���e���G�cv\��f5٦���M~�(��EY~�j�I=��5��// ��g����������Sz��Ȱ�@׃^,[���1�l�a����5t�����(RcOt��5=����*�W������vo�J���Ӽ=͐!�h }�w[�IZ"$����=�׸sD�zއO�э�+���a�-F�����ݮǴ��7�`����E����Ό�bqB~$������Y���T㽿f_���N��� ~�h�!rT2��Ur��A�'�`խe�]�^($����^�He�P�Р����@⊛��lM���}�2�B �
�o��d�Wc0�\�*31����M���#�G�0�<����G�%�@���bD�ڭ[8��pP��b�A���ޅy�eŊe�B�c3���8@��7W��x��2mZE�� �4pq[?�rFCX��h�����2�(v�����Wp�5��ğ�jX{���}����7.xX���a�|{�	���7|/�	����e���Dv�£aH^O,���ߑ���{�!�Dz�5+m����.ŷ�rm��F��,x�3��5AXK�x@��6�R�?E�Q��Q��GҪ^t�!_��4�x �d�f�s�����t�{�6/�q���>:1�U'|I��5�!2�� �#��Y(�$r'Mg��lf�
_�C�|в����ۏ1�K���B��0�4�h	g�Pt%x�1��{�N��9��/zM=�zMϳ2�aL�<mC��^T��8���1�b����Ձ����p�+���rG��R/���2)4h��	pA��Q�N�ɧ�su�t��m������3��ǫ�s���U���k#wI�r���.Fֈ
�շ�;:Ԇܣ-�3�ݞ����ߌ]�n�qɯ+%WxR���y���q����:�+\(�9w��eV�I4�B��7b漋E�T���F��|��X�c1X-��e`	!�7s��F6��]���.�K�����P��J��1ux��j�i����b�<ل��&��OO��R���cP(p-vc}#�:��Y/#�53�����sZ�=�dP���b#B(	�.��ˇY>�ߪ������*@LS���/`����6�L�p,��JY�T@ g��Q�iCk8�Դ!b{��jC`h�v� ��x,�X��^d�b�����.3��-p���������w�\�B�t��*���$�x,a�	�J|��5�������fQ���g[�n�j���V���\��R�!m݉V�(,wΞ�X��G��D�{��ƿ6qZ�\�L .�:��1KW�NB�x�8��{x<�U���PIv����>l!�L:�{#��E'V���ėAA���&���8vz��˧�Z����I~�/��
i;	^h-˿�f�P�
Y��E�|��r�#�����]��k�)Ul%��V��ڝm2}+��hb4j��SĬ�<{���Ą�t�-NW�N�H@"/ޘ��ǧu �Ƶ��$<�N7]��G{/8�� �K�FjSq=��4D�#�@6�2�b���ޜ�EW!�T[��ӟ���x�;+!
�� �fp�\���I�n{F�z���QD(j���Ak��� &����
��/����=���w����*�140���CJ���/
�:��yqRWX�l�|Xy>�i�
�ݍ���	��[H�ӈ��O�Rwo��%����"�A�R��zL�N#ȃ�6�)(v�Ni���qƩ��lw���v<l2>����=I�ű�(Om^�x�!�q#<��i٩F��DC|{d�@�C��ns-~c�%N8N|�&��k�ӻ�#�N�F�h�l�̋Qp��~�^�!d&�m7�,��Yb^���WT�D�C��s`y>�g�a���wU����z޾��"O�=���H',ɞѨ+�d?Ni/�2L�M$�vӤrF5��5�i�P�bbi3H�b8� (@��|0�կ]�0���z�r��F�WR'!s�=#ŵ�V1��" �Ve�WC��t�-&|�L�϶�h�@�\ D`͆L���K�۞��Vz�윾?�^���|��yҐ���#�wo�r��qR*g���'g�*�6&�4!k�@	�)Y��B�dѐ�v�F�S~�&G�O�����sX��0��W�F�]2APO�~h���n���*��jD
&í>;��5��:n��V��Uݬ��?��.��=����E��A����B�p:/`=�jP{r7�|�@��g��ĦY�hqA���A\f��N���D�]`m߀��^p�ep�L��A��:���'b��*�}��hx� �����u���'w '����|P1���=
JS�+��;�K="�g:(�2�v@����V��i$:�",�>���S��{�W�@<�����j)��#~!I䙽��c��4�r�̽�����G��OQu�y��pP|�*�KE��>�vh��]���	�V�!���?7��p��?�V ���d��leT�<����"�οN-�[���-. �Vx��Ҍ�����,��P����v�������l;�>è�
g�,�~~��%�E����WH������>_�+�hr�M�	����pAt�����<5ع�᳹���f�)\j&{��ؓx��O�o��"Uǡ5��X�VuZi ���t�mP̳���]������9��k�UJ4�ϑe�F]%��UfQ� �67��|^����f9
9�eF.h�l�����~��N�{Xm�&Sm0�>ɫg���S�3�Aڇ�i\�<<�]o�.C�x8��!�Km� �aя��i/�o����	gy
�1e�J��}�^'Ϧ�-yю���F��P!ǰQ��p�S�wM����f��}�3fW�\�������"���]���S%H����G��u�y�WT�ׯ�f�T��­1�N[V�+����`�Z&�������V^�)Ї���y��QԻ�r�t5�u-���M7+�n�OiB̾W�U��g	�	Op�n��T/[Y\���Hgr=.�<�a}�Y�R�T�tD��/�Vr[],��(����rdA@8�0�l/���*����g�h�1*�T���c�h�%��H�Ǳ0FJ����U��&%=��ك�8E����V�y7�}���V,�/��K6]cd�s y���0�*C��+�h�\��Z��R��98'�ܶ+ҁP��%D�X'&�-�/���X�z��ۈ���U��H���J�B][�n�z���rƧNX�Q��|��������{��~(�E$rƑ!�����q���p���CV�%(�[u��ح60;�ޯ%=���8~j�O/���4d�Q���/i_�8����2M^a��g1Vr����2S�]*�8X�Ŧ^�饭C�N< N#5�@񒅜��'��3JR����Q�,@Q50����0.�BLX�eTKbѶ�*i����F� u�z�J&*��-?@ଔOg:�<�#vZ�/�2�ѻ�B��ZQ<Vߚ�g���Y�'D�q��u���=1�|d�欛R���,;� ��~ǝ�M?0΃�T�xr���R�ט�l $P��fX�ny��|HU�o�9��-!�T@�tb��m�_�c��3g��bt|�y4 Z�7k�Rl. �B-�MZ'fajj|_5,�������U��(B��G�\���i��01�C���4�9��Ŧ��� !Օ�nlL�eZ�QH��P^��/�Ϻ��]W$�g��:�Cg0��3�U�+J~Ta^�g�*R%����N�bD&J�*-y���.:�l�����]ait9�#�;X�W/���bAT*4
��6�K����ʣoSb�`���I����	Q��!�Z��d�����߅������ �<!zr,z����]5~�(�ܝ�SS�lL�O[��qd��d�+.5����M=��wA��������.��U>)�Iz)��i���!�#nh��χ�BB��Y��r+���;��3*k@s�ca1��*���-�?o�R�Fg�S~b�W�z����{�U҅�W�҆����ى��� Q�����]��#���y%h�B,�TS#��d�����T4o�n��x/h����Y���	c+��:�Rc�ͅ�}RP��@��/������챹�Z��t�L*[1��M�#S*'Y
�Y�1=�G.R�}�+0�M�ӵ~�Ҕx�бc_�|�ɱ0���G	L1K��D 3&�I�q!K'l��O�5_����]���o����+0u���_�
��r*�>ȎX:b��	J�A�L&x�ht�n2�*d��#��c�C���O�ʾ�hq�^̰(A*�$������M;#��œ�T8s˲oX��|뀍F�Vs~0�;�� ��}�R�G����zp�`x_[^8�ϞJPq�|�5���(�;$<·�M0[y��C��̪��d	6��`̨]�5�<�Ecp�/<"�L�mĐKf@�S�_�"l����&!��R�S6AI�L��?�w�Z��Q�.� +��8#Q}�"�y~t�j��W �%���7 ^�O���=�«Sl���qb̟7�-D�`�p�:b'o��g,�6��/t����^b�o�t�G3�J%��QG[��J�&ȴ�;�cV?2�miz�?Ý���p��Y�����;��ą�$e.�	��EK��2+���۵�/E��BDE��YJ4᩼>B�ڻw�{FW��b����S�2W�0aD��C)��*�p�������!�� ��omM��+��pa񏒊b�A��2D�֒s��(�ygY�_k�%��I9��t	d�����V6{�K��,֯|�Ŋ�*[q<[��t����	=��y���8$����j,�Y��7�T/%^-�y{��	�Oʊ��.S�r��`��Of�%
\�}[�	I�g�7D���-�$����痭�=S����AM�����
j�X�%�bO�u'ۋ���������~JB�Fk�A�G��#pb�~�쉢��v?�m�UZ��_(ʥ�x��r	�xom��!-��ܩ|�>��\�גtA��)GK8�2���9C9��~,��1�'$���k�m�\��M0|�4�g
[=t�,��Iȏ�cG�Ĝ3b �f�Sk�<�PA�83Io���g>��N�s�p}�\x�7�)[.v�� ����H*5�kI�����;��ȏ=_���J~$�ο1~��g,`���AR���O���?�qG-Ų_eR w�֞;<�����3d,���&���������J/�fY=�z�ݹJ�0~�51?]���bU��Y��cXע�$$u}�I(�[�Q@`�uJ� �#rw��������rn,��h���`Rv-vO)�m�wT���׈����d����_�n�W*��*Ý�ߋӠNr˱S,DW��o�d:�(�\�WfO��L�hi~��/E��as�ws�A�;�<�+�u� Ǣ�� �P�D�ѫX���Q�- ����2���!�.
?�}�"
rC�;�@��?�S`�l������ߦPѹ|.H�75���p���r& ��`���L*ї<����,AP��:j�:�:�Om.�L�3��65͗���y8Hӻ^��'h��\~]�LW#����t
��|A,��F>%�V��$�Ӡ�u�F��vҍ�U%��yc ����hɈ+�r!g��Xcv(4��T0�jo&��pr��b��|S H �C� l`�@�R��?���8G5.���[�f�ʺ���zXo���t�Q�5���R���Re�\���e��z&GoFn���e������/1QCt3�`����@6�B�H�k+B���ԉ:j9d�������=E�+q������7g��%$����,�C�6\��xN�jj��3���F�'�4[��C]!�[��V�N����B�C��q���Z#���Iy��[�д4s'���%_٫��2�Df�+�[��5�ߢ]�=�DR�)�鴂i��-�jj�1���
������ɋ�����糅���RU)�|��i$z�]d4��|��ޝ��ˬ�����B���
�2>:Ų�rXB�[h�	J��w�+�:��.a���$�'c�)UA[*
0��%��F�EM3v3 :�z�{»����h��B<V�M��g� � �׬s��]��qM��,j�L���B�Nb��p]~[�����U�V0=�"�e���������v�k{	�q����{L��^1�m-e��#��ȳn9�!���Δ'����t�abiE�MK�5_�����y���N��/����9�t���(n�
f�D�Y���%��'���~�L�-��!��y�x�W5rv��R%?���fr��P�%vs�q�k}��~*�/E�h��s偦�6�/nUE��$1[����/�%���M<�FՌ��AuW�f*X�V���� ��TN.��l���k�4	:�Ec~ߪ8@!`8���\�$���|8:������V (�y㡭�4��/+�h�sXai[�*��5֍s��zezp ��7�o"�����fAi�����'fo~������WS0�J2�cp���ss��7�k�v�`#�
e=���O�Tz����%S�'u��겹X�>��L�we,��CffZiJ�AȶL�U�>'�mU��^��h�~7�?g��S�B.�1���dM}ZgDӕM�**  �+���=þPXXx+�_{��G��=����_#�vȠ���+Z�9Թ&R���b2��xY65�JM�J�<��Et>S%.(�!�R@�r"�����4��/�ׁ����Џ��{�7�ؘ!�`g�,<b��l̲��=0���J�w��q-Ųi� (i��Z��huj������a�Xb�b�ȏփ��dcɼ|Z��FO��i��ZÅEd�1�l�?�YF߈��#&5腍G�Y R�������e��)45��6?�N`�cLZocSM�V��EI�Q���!���P��?7�uA�k���ce ��[{!�)RګJ<remU����q$������>%=�k,��,ާ˚e1�j�3�����؉��H�U���G�#��d�V����/B���A3}�﨏�������,܋b���3x?<�@�V�lrN|�h!F�vv�𱆠�N�i}��� � ��ꖕ���g$q~������LW��pWU��i���#7�]M��� K�I�g$�b@�I+�ʹ�.�����8�<�������54����:؞hm�f�DA��k׶�PǤ:��?-��D���8ͼ}V
��uk���}Y$���W>&H��<efkS�Bo���O�'���7'���:K�L�+E����m�ALg�?��L^F��ؿ��F)���
/�����'��L��Wy�ƒ�1��,�	�i8	q�Tp�����,Vnc{���!��k�+Ŷ�		�}����+�`��BO�C�>�FB�;9#����]~mD!-w_1މ/�Q!*���*�Z����+�k%��H�ˮ?��W2N�k.$��wvD�O�"����TW ���VdS����Ƨ6av, ��:n��ln
QЈF��AE��q̵�r��W,��B�
�ZnT���V�K�Fܒ��k>M���*ܥs�w�4����f�&lN>��~����I���A �?#,���nTȃx �֢�zvs7(���Y��&<q�޳'x0�PZ)�l��ף����~^xQ�Pa񘬆`���r�}ij�e�ʼn
�N����.s��;7>E4�V�h�oH�i&]4�e��5ż�^����`�>
띍���1!C5�6�o,�=|Pz����*���_ĳN���=���J��uf-��H��p�Z��-��T�4B��1W�m,|Z5�Yme�'r���6	J[� �W/FԺ�qr@Ǧ�w�Ҭ��y���Gy�N]1����%1~��h���N����!����J��%��lSfP��I@/]_Kt� 2a������J��h!���f��#���^$OE�r�QA�����DL�蝪RS�k*��O��5r���
B!%ys�|\��/�F,L�C����~5��x٦�4�`6���v�-�ѩ��ÃBkxAc^�;GaM:2��t`�oN��)�(����5x1�0ďK��Õ&�ׇ�h��Na�4R�_�vF{�����]��֏"��]{YNT�����.*�H�x`�69�;,��(���d-��1�1�_��X� ]H��{;&]pp(В�h���H1�z_���W"o2~0ڴA^�M��&u��瑪z���{T_q��� ��^�ZΩS��@F�����,tsU��(����bZr�\�&��osrE��HxR���,�m_�gޑ�d���:���P�pF�Kh�Y�"���� I���V~���T1��{N��c����6��s=Z=��8�&툻uH�ҦCˍ�ܬ|�=���Ρ  t�#�����p�$�:i	���8�#�h��"����:�y���R��W�,=S�T}T�/8 �F�\b�Ns���HV����d�9xM�FbXt膔J)�C���~�����hyo#�%�V����w8�x�F����!�0@8���V �S���*'�fPJ50ᴳ��Z<�F�0(���U��j�-�씎/E��qN�ث�]�H����e��sa��]�;Y �R\�a�<M��ȓ!�;��n�%	���ub���I�����t\s�9}n1�4����~7�S ���d����P��غ|��?Q=)��G�>����-����m��ob�ӹ.a�La��4���~I|_�O 8k�t>��Oy�!7=}��Şa�=
��">�*5N�Q̓���J�^n�l���|���o���J�/���j�\���@p[#!
�!��E �-s7�N}ܭ��j'<u��9���+j�C�R�6qh�_I�Q������7����\,��$�-�ue�<�h� �",��ey�x�E#�W��=Y������D6��u�MB����=W��]���J��U��Rޟ^���R�! �A��qY��Ъ�#�m���T�
�+�@��U%V�°��ъ�_���A�M���f���t���f�IO�������?��oZ��b���'θ��"�)	&(��!w�E��.�$"������M{?�yk�C��3[��ߢ�x�͇�il�����K1H?��hv����}W�*		C;"��\_A�o�_l-w��7��idI�#6�����M?�r[�����]o�:-h;���K�t{oݭ��=8`%��تO$��8f�٫��q4�(
m �q3|��/p�,�R_�H��	�9�1G�D1#�e�D1�z$J�#6�cC	���Y�9��ICR�r^��Y&!Q3��u����Ք�YDD�n�"f�ښ�	��j�s&����0죊�"̩�CX�8fv���( �&p�Ƚ��(��w���@��B�O�\�NgW��rģ�_�-\�抐�g5K�r�_�n��{#��c7�Y��4y����k�}���� �,��y�[���+=T�s�WڽO:�H����rt��q�@<�_m���<_"�Y�J� ����(��纏AQ��-�ݕ�����\^#�f/&������Q��|kֱ��ǖ-�o2���<i�ђ�w�ȋT�7 /�V�`6��+���Qk�eH�z�r*Wф 
�����Z��w)}������W=�G
��Fr��7��T@`P9)F�W���v^�(��D�3NYd^
p��?)\������.S���<���v�X�V�9r��4Z�2&6�Uz�	����	*<���MA�[�/�Z&jv+�����d����$0[�%k����ژN)Թ�s���y��8{.x|�A6����$���bu�M��>��������Ţ� F�;�;�/�0�|��^)��&���*����L��s���8��~����D8#r��JzBr�n(�y��,�٥JּeEiP=4P�N����Aӵot� %.��M7vG���>.$�Y�^W��=�{Lh8J9�j�b�y��lq����H04� 3č������" 3�[FK�i��>q-t�+��@E�L��9�L&ݔ��؀��5dT`����>��!�A=6�ɹ��p�0�'�R`̀Q��`N�ǆ�	1NO��#�.��f��C���Q���a��c�@>�?G[6ӎ�ɥ����|%9&�����*���J�=� *���݅�)�JeV�^8} Cة�+q�C�jF�Q&$�F�O�4���ܾ�܄�cV����R���wPNA�bD깧� ��Pp8������s[���7V���=!��Pk.M���D<��̘�p�u�5��O�i��Y,$�V��|H�I���o��F�W�$*��޹&�z׾�e�1���{��q�����	�	I1t<��Vɏ;���q��(Y�#�t�\h3	=y3�	eG������P�O%1E������&9��}],����\�HPha×���j{?��"܂�s&���|�bk=w\�Ԑ�A4?��3ǳ�M=kl���n|������B����ˣ���ṫ�uw�5QNg%�z��9����Ïu�
̖��a�@0)*�7����(�~N��#�5�N9I�Da�Ӓ�9<�>H�w��pZ�Z-kƫh���ltt�@�5i	K!�~��������T5Z{T���ܨ��_��0�/�Y�&<���óF�`�Xy���8�t�a���<�ͩ�V{�DA��wl[��߇f� ���}�n �Yb ���Eq�O^�k���&Y��Z3���/Z�W<C|�[�����v�T�����v�K�h��+Oھ��ķ Z��1��p�)N�:��A"�b��C?�xXUW���zR$��J��Df�b[��Ţw޻�ݡ�I�\$&���PY�U�?��֒� !�p�8�nV^;96�eQ�2�1)�d팶��O��Ý��LC� Ev&��>2� 1���qF�zh.��_�]�q��H����,<�q��a���Cj�^�usMm�rPA�$�E*[ 3��"�?RL��B6��-�u�JJ�M���|���Z\��\� ��Mp�U�7����(�H����8�0r1�L�2k��ϲ�	�P����7�_��F�;qQ��F��6�Y1(e�C	4% ��`� F���2�;��!v{`��d��BdV?�tZ>�)���p)�FyJlZ�Y0�V����j@2��S+C���!�Rq��HS��v>]��$�ܣ��_,��tl���~�R��*k��ݢ,B:`���Q֛?V�>����^+�𢢩�9��U�?�X��g|l�m)�E�	�s8��o��.ԡX�J�b�=ጆE1���_�b�\1	'7���3"��ށQݟ�����I��/�?�z��lM�[� ��tg-�
2/�t�Շ܁�մ�	]��g���P,t5Q��Xh���ZJP�SR[*��8h�>�?s1`��p�yP��A��ļ�#�U�kS���i�2:��T��)�m��-���̿�3���_h���qۑۏ<-sݺ@��U$!�Oz�Y���_'��7�Mg<,�\�ނ���e#]��@�����#�t��&uP�����.�O�����[��|�~?
8o��&��n������?B��8��2K�<��B���L߀Ϳa������������7��(�j"qŤ�E��,�C �{iꡋ�p���̿L�ä��|:g��Xd�`�E� ��9�O���_�S�s�]K���`��� _�����<j�w�;cEN�;�1t�wQT~�ȮU����02�/K���9Į��UWp��=k�!�S,_���������J
�8Bʈ*J C��g�? �o:��;��V���n�}��]�C].�O�t�PZ�;��lu7d�M�0���^�B�����,ROЩ�rn`�Ϗ�p���Q�\���Lk]��m��ˇ�R��\ó+��#�`�i��Ӹ=kI-$��.[���<�5-U�6K�{�C��n��G���\�{ۢ'4�u�`��Jr��
��9��k?���.-�Im-�ɸ���ض���cJ�*l��%�FL����������u����].��3ζ���x��[^���M�Q�����}�ӂ�����(��4�ܯ��'cFCɾ��=��0}�������L�a_�u���V.����'pyp�kk^�7�!@�'^?Pח->Na��.f;��.E�kA�vd~[Sdu�Y���۸�<H�O��'�Ϻ�"�xm_������X#�z�+����8�R����oa��J59Q�y���-��IQ^���v¾'�]~.�D�LF�u�b͘���ӹ�@g��iF��L��6Z���:��RU���C��Zυ��귶|B�Y�����Yz���?�!��I�3XR���>Bl�wM�����x����*�~	��|�)�Io�vkA��$X���5��TÚ���¸�����C�� ��Ds�@d��3ӆ���놨��@�+)o�v:?l쭛֕5̞~~��o8'�}�I��bz�G)(�u�����P���[*�H��h��ӥ�vi��b1G�eVc�e�e�D{����9ZSAv��*p���2����X_vc#�|�F�6�|�������ъ���5,t �N?RD���a��z#eL�I�O�%�C�;�f	/��qش���R��,�Wt2>H���(�X�+��4'RM�V�܂T<@������4b��x��uD���<�T�0͍�����L���<�9�C�2X�x/^.��j�0��]ٝ���(���2h+h�ؼ�0/����W��|��Z�IG����s4S�����G'~�ƺ�[��j��#Y\��AtbC����]��A�c���s�3m̩$��`Ѓ��Q[�߈>����ߨ0Cܡ
�	W<T)�� � ����#"_��f��G�0��U`hm���)��v��c�|t�@�bpLu�{+����ьE�P:�+D}#�H��FF\�Қ�0	O:���T��a��(��)���C��U�Pn%�Lt�L1�|���l�Dq�1�o��W1��������e6�?�*<�DGLpl���r��/%+'�8-^)>hz`���Nu��2�3�.���6(HW��{P7���%��\ �L�]Gʳ^���k����y�5��G�	������O��E}�Y'�3z�3R�G� 1n��K�&�l����R]U �$q�Y2�a�Y����h�=�<����TGN���>�[b�쪪^�a�6��)�E.K,l�`����Y�]F�,�H*�:��OR�y��|�ϋ��prk��,�r���t���F�f���1��O;G��׷�9�ˮ�1+�uK&À��70ݓя��7?,p���]�N�"�N$��eB#�h1�ҭt��zr��v�o������^��A�F�sLwEG`d	`W��;��gq�q�"�~��\�ͩ\���@�§ =Q�Wl1�S����{m�j����bq��࣓W��l��+E��̯�;��޾R�XnnJ[�����m�s܍C�;����sޙܤ��G�ʲ��Gj3��,_�z�u���5�T��>ןZ,	�Xh��Y�CQK� G9��b)��,gm���5Fs�ój >�-!?���]>n;���ޕ��U)��҅����h&4��m�J�k�0 K9���bO��D/5��3���G܌�կ=�t;р��rX>�gW�Rߗ�֓P�
�SZ��>HS�c�&Q���'т*���/l0��h=������?3 �n�~v�����;��4v�IG�13�Z3��Xr�|�a��{���ke�Ǣ�Bd�[j�_[Ê@^�_�5�渙�@���,����!�Ҳ�m4�S����h�=M����L{��tv�XR��8�uN�طJz�h���Ϯ�~Y�����M�!&~y���NwSe�y�;��S�1R�p:��H�k���%�����z�����N]M�7�K����Q�������.����5���(y��͘��q�|�aŝ3�:�U���.:z�>����M9`SZ>r���XH������n�8�(��q���sThu!��������^�~޲J�b��)Z" �<�7��������B���Ɉ����@��d=��~4���hP�Z�uTx_f���e؊�����o����U{.��!�wMxj��<�~
/r�?^��i53T-C������Lm���<���3�V�zp�h]y�5��i�2o�� =��aM�ǐԏ*O&�G3� ,X���eLV�#{;�2W���7���e�^�J�Y�� Q�I]<���.G�MfN�ZV����~�8����A���ߵN@<<�f͟Y�9�4��vQ<w׀��X 5��'�����8`�S�����T!�m�J�q@e�(�����M����D��vȱ�r!'�Vy�}����NO_k��pб�b����#����\F�//�u�i�˶uA�V�k����ZAO����hQ�^O���W��<t��t�)ޑ����-�f=�Oh�1*\G���94J��Ά��c�3~JR�/�P	a��f �K�\[�"c��<z��t۱���X�"& m"���<j<O��ks��^H���C���:^y~v[s���8��h|5���ݍ/��Q��*�~N�RE>�����,+���6��1��B��_~��*�O>3.N�}N�'��F�Ǎ�]�2��V�Ds<��A_f�Ĥ��|~R&Lћ��u���`�.v0��%�d�Ʉ����������x��Mw�"�0^LލE��6Ϊ.[�e�;)�U��h*n<^$��J/�w|?Q���*�ir(4A�T�)J��YmK���L�<�]����{�8�_5ay��AN�'s,%um
He"
3=_�&���H��B
�x�}2����ZD�S�΄w�CF~n�ػ��𛾃W�H��<wgj.�*�t�Rm�8�3Ȼ3z����/�.��a-mb�����{�TR�>������R ��f�)M�a�x���|m�[Tx&�]��o��i�^��,�JF�2�����7>�c����Z��o����62�ww�Y����r$�g���q]�L�7�T��R��<c�%f禍4���<E����@����i�!�������ـ�seQ��d�Q�k�#;��2B>�*��������r}s�S�W�tVMH�0b֚K���A��@���`��tsѬ�]�l�I���5��H��ղ�#Ӿ%�4ӹ��4�f���Mך}�ղ���L�E��l?����J��߫25g��8��*L���/����q�T^�LGn��mf.d`К�zz����f��O�Q���w�Y��5�: 2t�4��o���m���10=;��F	CP|�	~Z�G��bۘ"�lwݐn왵O@�3��l� �*
�K�f�ޣ�+�� 3�="-r�9/g��c�s]�![�qi�Ο�E�G65�h���"X#�!覞\��G��} ȵc�px6𧼬9͌���֏�%>������K\��gٹ�h4\��)5^|\���`�T��0 F�1�9І��E%�3��y �NA�H��gR퍀�c�:����×ǜj�ŇdihA�\�VXz7[�s$A�����^Z�?EC���J��y�x70ֵ�J7y���%�J��r%��q�ޜcE�	�$╊��E��*���T=%! ����:�춞F��я �(}>4�0��'/.�⹁m4U&fCXx���㽩dćZ����\
�秊 �3G����d���q-k�婵��T����C�jt�$�"
�aX����-l\�ZjT=sW�i��+������]����c���?UC��s�>�ˋ�C#��zA}�ǒ�	�3���w	�
��jn�/g@���9"��1!>��a+�FZ���"���8;�W����څT9�6lJŰ-
��
���Y�
�'�lplR�a��ҥ��"6����Ц�&]���<�VM!o���9�urS`D<
`f�a̪�/EA�@I(��]:|�؝qQY���@E�%^����o����x����02v�(���������!�K�<��J�Lת�~vr�N�y�/��#��f��!���j:}�ɰ�)R��-�j_��`��0��Ί�$���#�(�L�~%���T�e:���?�,wT{jA*�����˺5t�&C�|��?��Mu�*<5P�� �O;N4�Dݲ�,K���?}�i�٨�Ϋ��1ƙzWK;� |��oX<�x�9��3��qF��AE���5nXM������{�ҥ� n�+�ѸNHMm`a}�a�w��	����.���ի��n/"��{�� ����'V���eM�A����t�4�T����g���Uc��oe[���
�Q�P�W}x���i.�#��q��k�#{�1�Ou�:Z�������9SC��&�'���!����r?��qs�	tj@���nu��H_����~�����,c%��)wt����>&k�Q��Y�8U#��XF���x��}�a���u*�͌��/��u�IDR�=]i�{J���
�%/eGӈ��iV����# �a`���
�,X�zv H�1j����铘RxJ*���T_���-��v5��e���Īȟ�iq��WҏT	b���N�,����D�(4����?mp���m�7:2�szZ�*�o2 g�������D�
�>�xo������,"�k�UJ0�����=_��p�����π���<���5X��j7���ؾbp��(ON,��Ɖ��������·4���1���Q��)y X=2���;����v�<���H�J�ڧ.�����?���qo�L��g��_�4$�dJ�O=!
��<q(�q�%m��=�׳Z+s�NȌ0ܴ�3#����T��d�?ʺ�Y{��юg�_�=]�j�|G�c\^ٶԥz�C$�/U��?�M_�`E)�İ����;;�UB�6�T1�GF�S���6�m�Ѝ\6��r���]�J�2@pL�y� ��xQy���,*d*���͊�; �7��T�m�o�Zs�Z���Z���"-����F�@�v4�"!�Gj���3���k.��p!�M��W� Ȕ����S�B��?B��������닂6�������j�� �?������Wp��@��&�%��t$�+��gตJ����L�:��2���/�T1Ț%ψ,m-�i���Lò!^�����a)���"�9Ko��C��EΰDo�����YeT0o�>��:u�y�8$�A��>�Z��m��@{[�"'�����^7��3������o�W����O��Z��P�ܑ"��o�%�&���Yfw�R�2s��5����v����I�2i2�[�\���=�_V�hNр]���[6�r��R����Ȱ�2�\4�&o�˦�DX�v�*�^�Y�3��$��%�"\�f9f����w�����P��#��h\�T^5��]���/&:J3t��9�Vb_3.��\^�6>'�����_j�U��&Ğ���:B�L2�8&��S"�.�ڗڼm;x��YsCd��d��$���$r�k�ʦ�0�SD��~�;n�r����v��,�ӽS��SuK���ܒ{�����D <�.l#D${+w'Rq�3M5�f.�R��F;�$��tK�D�R<1T���m�T�����8�ڮu.@<��t〨����ѧ��B���di�E)���$
��F8kq�{@?�~g:���}(
c�g���i�v��ðk�#w�m&SK�}��*B��"P%"W����Hj�/���JLԁ\
�J^�sr��JݷUf>Ћ>�p�B�~�+Ѩ���ՇX9�[�<|ͤK;�IjCU��n�,p�ih��|4$ᦷ\��M�9(���y�J4�aR����x��O|�F5�<�� �n�+'4��}�&�1F���G��7�߂���������aj��a�Z3[G���n�i�8ߊL1��*���yF���GC�1K��.~�
ԦP��w3vCdL=�8tH�|����%jX!����`wv�� �b�	�����+�W��٘��ֺ"�q��PE �6�j���<5�$���#�x�7F����<3C���}W6��Ҡe�&D�W�Cx�#�M~i|&ݩL�o]�X�*�C��=���Me%D ;�=i+��_�ǐ�cqI�m�^��M��6fXAq!�f3@�m�׾X�S��t�=�� ����U��A����`�CQ��b�j"p�ezGKkt��?��\1��UR�3������t7�����3C�/AN��'�B���Ȣ5�s�{3�Ǟ��P���jM�Kg
l�,91h���&@�_i��ou���[�x�	��แ�w�%�LJ��9�~>�س�	{`�E$a�K����h��yY�~�����O���4 ��(�]g��2���d��8�+�{�b�`�ZBv��'���o.�|PI����82�ߨP�%��^���ISt�vH����IE#�Q��ݿ�18��$�)4^�p7��,`f��x����-��'���k����z�2J�5���Nkf�bc8_�����)���@u�?_oiқC%։�4��E���	��!��\Z�')�?�E�RE�a��́ᙙVҁbI�Ocڞ���wj 6e���)Ź8cΆB�*��.�Ty���ӝ�U��F��Y�������>����c�(��3��q|ft��$������i���&��������Ԧ����@N����M+.@��%!�'>�~����h<�3 ��8.�eq�w=檈Ԩ�X:�R��	Qj���M)U��fR�?T�n\�WC�ȣF���m�4�D݃�?��O�h����<��y#��>�ҨH������'��l���_v����ϫ�����J�N���ro��	��P�[����6i#r]��Y��C�(�|-��z��330�J�m�@ ����k�m�ƺ�E��/S'�k��� ��(V�h%�����=���A=u2+w��T���n���d�rOH��^��q�&�e�j�~wuF�+�(@Q�Ÿ�Ӽ���k4ey��vH�v����3����) 1T�턹��Z�T�mD�޸�����/��p܂1�6������j��v�/ڱ?��Y���.uw���d_���#�j	%8�?�nJ�t"7à'��
�Xj�z��N��ˀ��7J���lct�����Bb?~q
�߹��}s_�%�w/��J0�}�D�\�����FI�/��r��N�&�f���y�;� /1nq!sf�a��1r���,��/|2Ts�6�s0v�$8�xT-q��Ar�c�˥/Ek!�� &�x}�+�G��`���܀����͓�c,��y[Ɔ3"��J�h���1�өIp�q��@�+����ŭ�qw�1� G���l�F�&��X��YZ�h���@F!���V�1����Z�օԈ����u#���Ҿ?�	�T��ͅ _?����H��u\�v-�7�- F</z y7\��R�V�zV��`a,s#�X)LT͐,�0��/��z7���(1~VY@k�k���M���	�Y��ZOT4Z]���
�g��d��k��<�^�8&�p /mX���>�䉲�rV�NƑ���РQ�7G�p���<K�E%1? �#�o������ ht�E��W�d��wr|xa(j�?!�x��t9���n�:�3�[���d���\R/><t�D�L��<
�ͰR���(/��'��syY�]_�`	{���Wc��|�{��F+f%$������b$
�߿7�&���[���ʹз�#<:�xK�����_���ݹ~L�	���MP��bR�Ok
Ls��V�4w+�x�|����IY�FO�����(���2�ن��/��}��p�`��� ����4���QW�`,�����CHpU��HxC��"��J-��E��E�s�PM�h��OF�@���G¾�Y�6�8Ӥ�6�p��%Jg/�*�����ƿZ�s�0���Is�j���y�`;[I��=Ҏ�Ux��sD�͖���
1��m��$�<dҀL$�?˅��'?J��2gla��
�ߞ�/��g�"��0�dT���n��8k첚��������ߟcQԨ����R���J7<_�Z�"=B���#6�Q�#uiV�mb߳:_�'@�q���ȵHwB��f�������9ƞ����k�IG6�]�_���k���)��I��r|�A'�^��Q�h�ܒ��bAn�}��z]��<�o�����_OM�/.�^�'��V��G-���x��wJ��Ǆ,����V$��Jz������#p��'�y+�e5mMq��sA%�d&�'������9��w}Kؐ������@�{��s���8t�$����n��k|�٪4F�ء3ג���3S�i�|�Y
�7t��z2��,���>Sͷ��v5k |#�a���ܣ�/W�QG���L<�ܤ��TK]�|W`��Y������mb�?�pҕ�4�D/ɠ|��Ec��O�gu��H��86]y/�;����6��	7"���1�N�G���U���A��k�>��'�mF�9���0����<�Yly����K��U��3�O1�ϫ����BtZ�/Zb�d�B� Z�I9�ps���ՖV��i���n:B8����启�s��<��(!����<"_@�M+�}i��,�nݬ�	���W��%��Fؕ��+!׭[3�S����Ԧ�e�hf$��<�g�b�W}LWea,u<M���,צ���*�;G��8[}Eh��O�H�;43''���t3p�W�2�CO��J�50oz~�j,��t�M���81C��S�:�o�
'�{=���L����my5Ԕh�GL�ش�^~M�;��؏��X�.�x4�9ۉ�l���}����M��ߤ�!f�`����t��/��ؐ�j��e� �k5���Eh����(J�@�B�wW�b�r��p�>2�
ݹd�����?�ڮ�y36� `	��9�7oݫ�ڞ�{m���7k�ta�9Lk��I�b� �����PG!V�
.�K�Y��7H�Њ�)�̯�k^A�%`�X�ƻb���<E�=��}j�6�@��	���I�,+Xng�ɨ���.t��ƞT�y0n'��E���R##2����L{p|�0(���p<2AB����:�55�
�L�����qS��u���Gu^<��44S���<�{:Y�/ק���U�	h��2�y���P����o�:�ͦ�5I�m������P���/ݤ�]��qn�')��|pO\6�_
�UMC;���R1�9u���+b����0Jpw�@K�=~��=�r��57�����7�o�9ڒ7Y��Qf���������<��?���k)w�-;r=7�*|.�E&�dx�pt%�<hs��m���:f�Z��/����5�����=}-^P��&�T�:S\;�x��t��UA���ga�=97��E_$��r��]��Fyw�1s�!X���Ȁo�URRԺ��Q�r�4ڃf;@���H�E�N�w�ϧ-w'G��þ��d��o�-�Lw���It��U{��:��c�H��31��a�򊞤-����z�q~�>C�Mp:G@7ܙQ/SJ�6F���������1��+�a�Щ�`1>�5�K���9�#Fg�|���צ�k�0�S%��''a_�b�4��)IC#" ��*��Ћ�T���ё�H��?�W�]U�?1%ʕ ��x^얶9[bND$|�O��5��Y�<2�Y1�J?�Rg{G���_:�N`�]R���;V�����I�tk�e�Ùٗc��xI�hu�����������_b���+�-�����z�A}e�T��w�����j�Q�ɋr�����_��kG��։���p�93%d�ԇ%H���.wr�{9'����xN�vξ�w�"���Z�H</t�mP��5w��M�V��o��䚪Ls��
<x�t�I��5�v�	�{x��OK�J1��<Ca����Ĉ��ip��8��Uj��7;6e�G���wv��[�i̌�7l"�Z�Yiڗ~����W��Bsѥ���;��qLa��stʚ�)!q��z�Um�9��ҡÚ���G�{�?�]�� w+�[-	0B�F��e1��q��h�))������g�P��d8��um���R��_d��w�2d\�§� _pet���J��Ƀ7%���ߢ��-%f�@ �ʒw�����qvL�*3�aM���&�C;,�|5�t�O�����K����KU�b��iy"~�U�j� /���w��YϽ�IB��P�hV{K�ݸE-��]���>�+��������_��ydZ�3>8�Sv�R8��r�J����[�J�.�چ�V��zY��{wguNb�x�o\e$-�?�A,/���u��,�+<��
�� �o�[��:>���ڄ�K��#t>���P�d㕸d�@*4���E*Χ�Q1bl�8c�ɫ�H5�I\���;���=Rݼ�y���1yN���/iX�0v,_�q�M��=�l�M�O���0����o��~��F��_�����Q���������ؚt��2�i�|l�')f�p��t��d�f�37k`	�r�<4!�áF��>����	��S��0X��:��y��'��JL�uׁ�����K���E��v�ܧI*;�����J-],QIiO�&1��A(��T'0A�k��&���m&y�̙d�����U��f��-�w_�G �n����;iy;nQ�x�t���5*��V\[R��$W�x��JY�;w#/&�%1���k�)�5@�q���Z�oo�O���~�#H��t�������&�qYy�T��p貴�Qnc�ҕIQӑ�����ȿEt��E�e��,�"�P��<h�R�Y�l�gvp�e�ko|^���ɱ�j��/x��洓W�ŭ���[�N�N���'�Ӂ���*Ml�u�FB��Jr�R�uB�d}W������-�����ڨ��eF�t��f]|f̓�+�D��g������ڝ��Z�U��b>��Rc��٩��ЋSc	 Y������Su�lv���X!�(�~��ͼƁ�2P%o�7˂i�c:`�C��z7�C;�vY���Ƞw�舛�V��[$u��Ԅ4#^����26���0�� �O�M��@HB��L��bJ�~�g���ok��t,r��c[՝%�d�]�,S@zP�8"��n�W�j�3(�ڳ�ʒ+#��L�M�F�G� ���y	t�^ACQ�'u��7��R.nEg�n��tL*�}t|��:©��G�'���*ݎ���uo�|I<�)d�i�D�Emb/�csZ� i�>�c�d;�1_9�?Χ$e�f�(�Ch�1�eȝ��
kɆ�M#�� Y���~���T_0�H�r���� ;S��K`��B�B�Ȥ�)���3j�%�F�� �Oi)s<w���5�.�\_x�ٞ�h!�
ơ��|#/To5��7W�k�Y�R��C���N"�\㺇����j��9|�;�5V�r�6���P�c�q����>�}H␍+Yw
RIj��{�!'�yM)�W�i�1�}AT[�cv��ȇ���85$˪e���>M�;)C���!��j�?8_�Eo����m���0t�����^���l��,�6+:Z�,<��oʌE�PaeQ�����Ϝn!��$������1Ѡ����|�&�ͨ������J~�w��.[��j�����)��0JL��0�p��'�[N�Q��a]�c0U��SL4��fU�ʫ1I2�$?פtf=���w��6FL �e$)��̍�K�3�|uʡ	鷮�[�?���������VW�e�4w��:�\��=�)O`�1�Y՜{�@`�H� p7�>���Aw�D?K�b�}~�X�s ���0M�p�3�x�(��ӽ޸nߔ;+����[K0�#U~Jh�`Ԏ���K���{#���C����5��PVX�ĿZ!d֝\����E�k�It1:���W-{SQ! ��k��yE� B����p�����E��}�|q��0{�̍���w�E�h���ug's�۽C�4��?��Ef���c �aT���J����ѥ}�I'��t�MRL�g��~2�E�1���vyU	ʦ��o1�����p
��`I|Bu�=��:E*T��4�H�p�4��i.�t�Ҵ��o ��ģ�K��;�������S�U^Ue�ؓ%+�����3s5gM�%"OD���V ������BP�R!Y =4t'�ڏ�ɐ�)Ո��@a�u,�?�!]�0�e��1�����\-������z��r����HI�f�a=d+1W�MG�$�ME�/�c����`)o�b��Hw��;I�?�S�a%����g.��@R��*�^@��N�8�Y�
pIh4��d:���GS�y���5��
�!p��42���o��_}�f�����I�~��oU��efS��q��Q������V���@�rW����I'ewn���0w�2�Mnm������-�Be�O���6?�Z�4w�F��C��[T}�H�]Vm5#��4�:V�x�e�{��� L6<��/Ț�L%�J�x�"(�M�[I鱣@��W 庉�����ѓ�9Y�n��aX�c*ka�]���<�ڄ;������������Q��3(;P��] �h�[2�(
���]��~�X{�p����X�'ͤt'���Z�{�F��1����'�FR5���~[����|PW<gFדUE������I���R7�5�ݐ+H��؊��/������8Nb��˪r��h��NK0��J� p�ts�� *z�Ul�I(�_/��󋷃ث�&V����:��	".��`�#X�C/�u.�h�Y�E�ì���R/���6'�y��ȺPҩ�h|�T����%,��
)��X�a+���ܓ�� Vͨ\�Y��2wD~�U���M&�}D�f69���0g�8#�X���>q_��gg�Qr{4�9�?�>���Md-&2�S���H�L� 㺢PhL�@�q��+�-Y�;��k���%dP �����������P����v
����`�z�9U�U��1`�3���0��Ԉ�XPT���F�k3!�}�L�;϶E����G�� �o[s�o�DQ�<���s��M}��I�����8ȹ�R*}��PoY��870�Ɩ�g��u���b3bkC�#���c:�c?�iT9~�\䪪�eܓ�w�ZQ�������E�IWx�a�ԉ���3.!���@:)�G��	y���:km��t���VcA5��+�ʽ���Z���Mr}�3c���� 5�����B�B���1��Dbԗ�X0�� ����a���s��j"\]��ٳf��~��=��*kAo���5����,
�J�t'��E��5+-��p�z?M���c�b������A�+\:�����I7��˻���H��"�l=���.�@ص�8iB��J#����r���p���J^UO\B�f��k5�A9�������o[纒@e
��8�7<B�g��V񷡪�[UF
�m��kξ�5�V�At9o�8�j�T�e�a1Y����e�"���$F�|IFv�T�'X֞��]��;_i�G����J0�|?FS�Pq$(�^�P]<��&�ɾ��6�Ӡ���~l�kV�Q��"�����i�s�_� �ː�r
�n�o �e_=��G?�$MH�8�TO+|&�	�w#dw�j%�W)3i�ͭK�"�d8����I�����PI��<��4��?�k&[����)��	P`7~��	����ysFH�F��?Ʌ��qW�����3r��������>�f�o�+7�B�A���~ �?�ʨȝ�lN�hGr�`$_��&�MDr��Z���.�Id����m�͎Kp�h�؁?���!�}��<l
+�l�fB�&��Z���3�ژ%.я�mb`
H����ѧsG!�	14Yey5����.Յ b�h���g$!�
�ﱴEd����mq\�Ģ��<G�X@���z�[���sXz)�B���S�������g�T�'v?BS�X�fU�y�܀P��l��bR&LO�/2�)0!O7>8��(O���а�1\��:r#aO�y�f��`�U�s����>P�O/�Ӹn��nW�[P���j����] �B��}�d3`L��B2�&YV��x��(`a��w'*r�\�"���b��}N��@��o�tR��?|�� �"���u��H�=�>�G�6+�<�^���n�;���bҌG�� bP��/G+���)?�\ݸ�.aM��95����
����tk��ӿFH]g�)ٰ>����v�����d�B{����Kf��}�F�'8"�Q��FY��U���,�p~��@rɆ�7g|���`<q��wO�U�m� �W��>�jPmk΅��D���Z<�����Q��)��2����n���v ����!�$��a�ʮ\��oo{63V�J��g\����x�b�6�ePTDd�S@�����в�~��(N`0i�x��V�����	���B�n|@��¦�+��z�w�81��@�s��l�b�q?�з�����%�=��Y�#[���8_��T��YwUp�/����%m��]��;�V�}?i�K!�|ZT��2)z�!�/_̀�<�DV�?$-�M瘀�C�&��D���Hn�6�l���>KbO2����9mU�>v�~'3-{9��F{{��)�fW��F�$D�o����y�dL��s;A���#q57�!���	S ��I�)H��
%&�
��WH^��^	�_�I}�H`3.���=EP@�!u���༔n��P�O�ݻĀ-6Ŋ���|�ń,�@'�}��co�(�:G�)h��!%I��1�C��P�D��lP����\��g3��~�L��r��I���o���*��}��l�+�u���1�t�+��������<'��P;�"jO�5K갵�Щ�<FX���g#��: [0��L!��_
b�T%$�D�[9�/2ff{�����CM7ǪŊ[C�'n=1�����(qr�1���-���L�Ĩ�]��G�̖�a��w�Λ���e���ow_�W�~q��2.i�#��5ܾ���0�m����=1�x��g�0�(�Ȗ��̥����`�ZB�9z�� ���
:R"�M�\R�W�c����e13����_#�R���c#��{E:Z�X���30��~��Ъ'F�-rOAWm�E��>�BL�.�VpW��1� �&i��f<�<Ye��$@��p�'w��)p]�`v#��]\�1�˂��2���͐2+��H�����{���u�cu��qdGq���>��Y��l��xlE�p��%Ae3�e*!ao>��(�9��7�Ɔ>��2�0hL�-����Ő��@9aX�0 �Ӆp*����ԦD���,�ң~���iذ�*�9��8f�}^x�5	Hn����MV���<�z�x�N\W��H�� ���-gMy��N�3J�����S�,�d73Z��F�{;�z��E�����y#Q���Uh˯xT�WS�
I��䓉�@=gWs$���'}[^�=:������"��,�̄�i�\[�+�O��y\z�ӻp�Πìb)9�ݝ�V �����5d틖�}�ܱk��ټ~�Ck�g�V�L��Fbhٖ?w� 
��t��U���!���R�(:���A$l6q�W�L�TNĄ4�-&i �8��WC�*�IRtTl�"0	e��{2��K�����]�m��+�p���2��n�_����Q�o�����6G+���!��!3{4��+}�pL����[��Nj��#a�[a�c�W���fx�:�o�����Q>�J*Z��i�)�_6�H�\�\W�Ew��˴��7u�=��lg�;��{�˳e���,a�>���i�V�8tqF��Q}/xv��	�;��C4�`�x���SK�-
BW���P�j3�P�I�'B��-�v�;��k�.��r��ہ.�1��LL�B�6h}�=������Z�a����ޞ��	~/T�q�xۑ[�v�j��kߵXWb���t��3x�m��[��2�Npz��b%�����xd�T� JX�c�0�4q�m�G^�8�7�oxx*���+9*j-y�P[�W�x�3V���hNC�0,d[&ncL��:�~�|*����b�� +�wB�꺲V�]���r�}�r�l��Άĺ樊����%*O$�*X#�K=���?힝2!&g��	�fky��8���̾��Y_�J�n�'l���姹.͍9�><e�e���U��-�"�90Y7��-�-�Z����X�:˳n�!�� �77(J{��Ԛ�|����1`�>+�Ss6ZQ�j<(.��;OӇ���[�6Ϝ~��I��	PW�os� 2�8�V�YL->�>��k���1:$��\�78�k!>��;�
��T3�%�����97�����m���~�FY+]yo��2�V D����T����tԡ����.��y?Lq� �w���p����~��c8D��tٛ�k��qDp���03K����ʭt��*���~e|���AJ7eUd���=�-W}�%
�ӭ�Y?+���"pg,dv'g�댮���F����=4P�C�
�@>h�k5w���(��#���Zu��(�f��1�FU��Ѧ����uC�)I��ad
�H��yd(�׭��#�0SDCt����_�̳z �w���J��Ơ\Gʬ��M8�#4�����R�R���Q?@b"Cd�<Lj"I��a�Gc.c3K D�7�#nu)H��0m,�|�X�h�� �[xE��/֭i
�EqOQ}�WV�l�<�QXR�K�(Ѐ��-���.���"�_���a��h��8��R�T]5t�/x�k��Z�B��g{ͭ��E{���O"�L���`�J@M׈9)B�W3��S���Lm�>�� �#���T�
�*i 1i�e>��*>�U ش&5�[�#\#	�Ms�w"zB���O��D�n���l �O�Օ*Ëw�ǐ@��?��0nZ�{-�k�Do�U	6�%hJw!ń�/���I��կ���v�z�Ej���i/�����b��`��D�\�90KD`�h�uoG�s��������ʮ�o���w+緂���x��yJt�,U�O�5rB��*��0�u뱜cpϬ��ރ`���h�'Q(��T�T�{��$F^���~�TN�������1o.e ��/:�7�o��ˇA�D�y�2�^%l�B�k78�Gg��b㳴�d�W+�%��Tn�wWK�iLK�vڃ�<ʔ�3�>�u/^mD��~�2���a�����eK4����ǌC]~��L6��֓{���'�������y��wum��yGi� .˯l�nV��g�:�y���>�d$��>.�����5V�L��J�ؘ.��e�o*U��@�/�~�/�˟�-������	��*#��c^wh�]�8��0��d)kYC8��#.�r���M��{^��H�?�sF��*tv���Z��ّc������#�ֲaZ��=3� BLH%�3!�[�U]@�S�V���O[5�=�Ũt\L��=�T�K��2l/g��x\T�
��k��N�l�Ǣ:\A9M~o=��u�S��u�\���@��_����K�X�?�#>���.`���6E/?��{��������]�c�9Q�)ä\��rj����3a�����MXi����km�5�[�\�oUqZ�'P���gf��m{�N�;�'�<;�G����F�4��{w�i:�j��0~� �Lܴ���D��nK82[���ρ�z��i�J�M(/+
mN��j�+I�*�4�A�-���p^�:~]��zg��l��oG��>sW4 ����ꖡ�s��A��5�Q�fbl�b��)��DPK��o�Ӯ�~��Zlg���8I�]wQ<��G�h���prigc�$�!T!Җ�m���d���(�?���#�3uy�mڶ��ٶ+�@��gy0R��^ɵ)�z[n~)K�T�V�kKFZ�כWmP�V�*W*���g�H�,��+�E�����8.5UI˔�H �LL&V�)qa��� �n����V#{j�v���+�Ǳ��-X�C���[��{�}!R���ӁjܚAZk��	�I��{���}�d���1��l�=�>l�g@m�Sk�~.۽w�+ 8�KD�t~`�8��]6�K��.���& �ef�CxI��u&�Ѳ^v��6S6e{�G�k�/DXu�>i,�Y� 9k��\^��m�k-����߮��cTf�#@f���Dը�P\5���Y{H˟�-a����"�f�4�sǅQ��#���~��37���ta���1>l~j�)=X�5σp�s�NǏc������2pk�Q�y���9c�ꏇ���G��'�����#!��ض�z�w�(�	j�j��o �I�/,m+z��,+���tV'�-J��hk�K��h�Qf��2a��04P>[�Wl�G�zxd������{��j`1bFF�*��W��x� �V:���xŋ݀�lv��?��FO�6%�����j��fF�ZG��9M�
�+;E��{.q6=���y�,��4��:w�g�_p)�Lf#�9��	&ˢS*���8`�s�#ϡ�����"�3m��D�{�=-����]uy��O=v�K^LAس�L���!��VaeLHf0T���K��t��Q)PSܲ��m¢t@�go�,`�	�v9��	K�pI|m����D�
�0�c�3�b������ØL�b�q�7ɓ~=�Mq'�SiU�ǡ ��s���?�a�}��^ZÂ�/�vb_UA1�Ia�#3y?xB�49�Ni?���nh�.&p��,�4rP���t��n�
�I�(]��%�լBM5.HGb�_�.�XQG����rb{C�}�-���Ԗm}%Gw���%���j�X�8���0��pI ��,{۔� �?*�����"96D�����7�8`��q�wI�
D�{�w�ei�5u)�V�8�D��$UA�0-��/����@��!��m���-���e�����,�&Ch�iv�ƄK�i�mH4+iM�o�"� oG�����Zp*«��IJ�	"�6��ޚ��N���(���ј k������;ta��W-�y���*�.�[��Y���0����m����E�ݴ� �|�`�$�1�YǴ ��Fe@	<��S��Ɇ(�uFWR�:tA����sc�o1h�6�M4o
Zm����e�1�*{��4�Y�ї�|ZK?�T�v#�m}ߧ����Uv;{��xÛoGC>�E����a��2mt�ۧ�H̉���d)�N��2-�D���g��,1������8���J��Ui���\��7�V/�֏�&L��9�'��J�?-�5�<�H�i��J��
(�b_R��#&���f��k�b��U��u',ʄ+
�0G���Y�j�|X�����m֥�mr�r�o/<�-@8�гgS9�Á��%%���U�[��]�T=3�����U� �'��
��3�룉zs7������g��
���%�S^���+��t%]S�����y�YR��o����=�IZ�����K/����?K(D���8^É̬�e5"��]+wh~�f����0Y�6O��;%G;=�H�ܼOY���ఛ�a�I�r�`V{Dz��P���*`��O7􁦼�Ë����&�+�뀢���wճK�Μ��1|��s���':$����O�W��E���P����]S-����WKR7�3��%�	2C�F��Β�Z6 �B�MA-��3�l���4��[����X�1�<n�h�u0B�n�����o�O�,�/q&�5	q���[�+� ��Z�jt����J�^ы��< v�,f���}�?��UqMx��Q�̺�Ǿ�p�K�50N�e�?	��ݧ�O	�4�J�S�1�T��q��X�qkտ��M���2zk"-�\�.�����v05NW�*���������u�c����pj�H�T�9�Ϫ�m?��={yH���|t�dT�{i�L�܈�x�}Y�K��.x�G��Ƶ�v�����"�0 	}I��l)*{8)�� �LB\�~�˾w����Ȯ����/0�@���J�}lE�p�>�����V#{��	a��^D�s���+DZ�o�w�����I�V8��HWa�j�my)Ȓ����������.@�)ѽ��?�ʮ3��e�3L�N���d�ѡE�Nƶ���^����3�3_�����(`}dZ� ��:@R�v�|U)5� P�C�%K��+@�3�I��v}��J�dç��(Ug�@�����S�%�2d�x�Ή��~̀�5M�'i%���~�{�'�Ώ0A5NXz�����[ �����R��!^C+y��ժ�nrȉ"y&9�����]Cz֞���v�E-6�]�W��B$_Wy�-�N_�I��S{�~�#c\�����A�Mn���x�-�5��~0���7��6mSq�UA��=��gMR�3�U�b���`s�Y�-0���u�)/�qu�q8�e�K�~aV&�A�.�t�$suNY�0\X�^����	����}ct�X��!�,ս�z4^��k�K\Ec�g6�"-��&��":g�Z��R��a�����c�������rw�ڂ.�gtp��7�J�m�}��]�ǘT�@�Nx��PIױ�M/?�R�$� �b�b<-���h�$$�n`q�+p��"J6� �.`��Æ�	�I2��}�2�L���E�	���ݰ��PX��T$�\x')hC�A�˩ߝulN}���.�L����J��w���4��$X�kR겂�.қ�Ӹ�9��:)�J�F��0��D�<㧮���?!-r��6؟��2va�7o���amK;dw�=�,d<�. ��CR���p�#���H�D�ż���(�q)θ��Q6O�V�����q���')~~(ԍ�v�
�>KH�BD�
G\O�"�S�K����JӍ`��Dω�чRa��y�8�Md�3�8x���>��>��!!��Y�x&�r��"�hN!o
���L��o���B%9�W<�����$t�6����Ȏ����i�����yMC���pO��$��1{O%E��qx��?���{ѭ�cK~�g�S�۠���x�oB��n���XL���%^���������-��C�ι�l��k2-�Ur'9�A�1�{�gH���������������qU�%=5p�%4l�{�nh�j�����U����gǼے47��,pe�>���)ҞNn��
}�!����G�R��Q<��9�'v�����T%u��p�
>����I�vN�d�c��)������.5_���N2�ɣ\G3zh�5����ܞ�F���yT��Q�I
�L��䙂1h��r�X�[:Tú$�ɹ~�u�ͭ�,���JY�\�B��Uz��j:�߬��}�m$<q��sx�S�����t�1Em�jy������k�4<�mVMqN��Ô�'p>G�@�
��b�	_O�;i\`�$D�kq^PuE-�S]�3���8#�ټ{�Ac�g5�e8�����3�D;������X²�����	&�m�~���	l)���8�~�!*�p��2�qCv�1ܳ�).'�r���:�A��@�{�jt7�R��GA��J����w�ۣ������o3��%�ѹ���o��GKܠ�s�����!�� ��J�SC�7�/������Î����.���;1pS�In�
����CcxA���G����E��B=��Nҥ�*D������wөb����i:*9����ݰ���
F���)��48I��r��' ,��>H� s,\�W��Ց��ZNi2)��=�H��!�a��B�҃�hk2�
z��w�C(S�y�Y�
��A=HJ�Q���^�`�u���HO�-��|��1xe��߃A����*�z�+�+'3����.��dq�*_@4���%4����BK��f�U����V�$?^U��@�{��4J֦!�2%���m�Q���\e��w�e���h�副-��WM�B���-'�H-�Ù�P}х��I��s
l�\$-�[뀇�sE�(3���I2삒���A	]���E����Ƥ/eW�4���a�=�n���m�=� -H���H��T�d�>�l�����P��05�#��`��í���a@��>p����Y�\2�#3Q^��8C�г)B.���/�<�\z�ޔ+�]��q:���Uh�j��CqZh{7!�z�l�(z���1�f)�?B3E}O�M7��o8��l+:��0����F�*#<�����vk=�N	i2�t{Ю�!\�
�C�HO��@�M��<�+�M˲|m���Z�X�MӚQ���~��Z�<Z��f]�б�G�
�3�L�Ì���RC�WN�I�4
�a�v���7"8S�mt� B�uq���%��Ĝ�㩥�qO#)�2Vͧ�sQ�L:*�R���l9ds*����#m��e��TР4#�H�|}.�[G�^�0�G� ��*$�`Nn�hn��	��xSG��ׯ",U+��d���1�Nŋ������:Q
7R����]��q�1�J�>�-e'A!H_�,s�'��9��c���Z1�G8��X��;�xM���z�;��t��	�Ɏ�ѵ�i��`�o�B�^���}�v�������è�Q�i��z��l@&���<�Y����\��c�'o�3� �] Kl�E��?43?�Cv��DW#]ը�{�v��u��+��>ّ.C9p!��}��wlT�qA�Q�~���D�\�C+�F��"sj�Oѣ�,R�3���䘴��AK���|����oiӘ.^a~������IẢ�-�b6aM<�z:������K�@�Y�X =u��n^$�NL$��:�I�����[�{1h�?T|��\`�z��7�b#j�D�u��m��J%����3��u �;hZR�D]͎����F�sf3}�	^��~�;-���ql�rhf���ef�q�G����g��T��5p����n�Xs��`s������*��钿�Aˁ~���=?��?�������8�тsM��Z����Q7������0,C~���U��	��4���-G����ur�bz(��e�4�.$'�|�҇f�],d�AmYjEN]�mx�i;���؝�PW�ꀣ��ⷬTo�/�q��S�V�w�l+��jV�ֺ��󷯳��/�k%�����߇�s�]$8��{�қ_�?��O¢�� 	��;u@KPFJ�~�6�EL�sJ�Hb�z���`w�z{�2[%�bp�&1�;��7Ҫ�}���80* �FL�3�0 ���.�>�^�"�7�$�zT��B]��
���{�Pm���ϯ��K�bm_���j+#�C�ým�i.R]�pU�HS�S���M�W:~��>�p2:�'h��Wǧ|ԟH�/�Ɓ�%\2a$	���.�.��IuT�����N�@��R�Zv1j�xfgʸ7H\��� �M[6��
��v>�]6��E��=Y��Lw�����-7y|�n���'��Ƿ
����HX\RŴ��p�-1�_N?Y��=�ٍ���1w,-��TK��Vw�#�M'��DcI��n���;
�B��mC����Wa����j���_2<J�A���z��:��UGฒf�)�I��M^H�-��Fq:Z���[S�� K�l=8j6OޜeR�:��Gg�r���>Ƭ"a�S�ph��.x��4�n��@�@�84>|�U0��&�D�yo�jϼ[���R��O��J�T��>h[RuT����H�~JJ��ҋ �vM�'���omЕS_�����O��0��4���8���y�y.)2v�!���DR��p�@#��;e�.� ��V�ɠwh�h���F��)��!��%J��w�XǸ�E]����p�N�˩�.��I�N��N��-ڹ���u2�:A]ɏg7氩��4�% ��*��aF�M�'l���Q@�QQ�T��	�V�sݫ�1�r���K��S��6�9�	��q'�`����`%�i�p̏$�'����C)0�*��S9p�2K_��[���CW�P��a@;��w��Kq҈�;�5��B�2tp���Ȑ�5����Ҹc��{�"[�H��Z��J������E=�X�\\��#9��>�T�'hn�~�W���Yn|y�zI�� �8�l?k��n��k$E�[3)��rO�|�]�i����J�����b�<?���r	���v�1�������`r��s���Ep�P���&��ş�C�.܈,�o�v�Db�U9j,��QP�m\/��V�ް�^k"���^S�:�Mm���l)6ȟ]�w8�ھ	.�+�!�3Ҡ_�=F��&�|�k2_������m�����i�2�����C�$����>�6m1/�<ꆷ���W�s�x��%���Äd砲�	�fۊnY�����A�����hc˒���X�-�Ǎu^��_S(x`A��ݷ����\`�ک{��Q�8Ӌ�6O���`�z�aN��@z������(�:�ZT�
`7�Fo_.�Q)Yj��K��N��6F�����p�)��l����{mKf��VJ��l�ĝ��V�8C��R�	Jo���X������e!�"R�3�֯Ƣ���7����{<mc����}�!Ev�<�o]���[���X �"�*��i�����j��WlG�+����u��gO�?w(��,���l�Wvu�c��J���,�^*�4)=�T��Ę@� ���Ǫ�'B�2�S����D��[a��&+�4^�Ɨ��%ګ���$�tl	��|eIouߠw,幦܋�R	�Q�4�w��R�Gx����']�Hu�<۔ѣI���&/`	FM*_��5nRF
Qa�?Y�2�8��a��D��"�G���!剂�<Γ�L]7E�Խ;�7,�"�y�� x����`#ǌ��_�
/�ViĽ,t��{ø��^�G��e��q���sJ��c�Bc>&����Oy`�H�n��FC��J=JYX2$�P˔D�S�$=�&#u<��P���&���+���x3*��i�_�ٺ�6b�Sb��#f(��D.�6��G���Ԙ����/�e�1�
���tP ����8#��L|:�1�a��M�J��Bn�ȣ[6�m�>Q���,'yl�ȥNmn��]�M�E8�G�5,�h���<Î�����2���ii	K����ܛ���R�r#��E�f2��
]�yy0��R��0h�p�7F/��>i�_4��d�������B'AE�f�z D�Jx	�������9��"2�Ü�� ��7�G[�<Ѹa��`��m��!��	������@Q&��.�#h�ר��؅:��!�z%�hr�qd�X��q����{SO�H������1�b!������躇���V��Q����=!R��W�T۝��Y��ک1-��xF�{�B��U���"c�����9*��1�yQ�=���/�+v(�Ie�%��N{P��`��ݬ;��N��;�'��f�Z8[/�&\q߶��6f�荽E�+����W;y�5ejp�%$A#�|uޗ�@�>���"� k�N�5aL���U&0����B��@
U���� ��]�}s��/с�@�7����-
4qhpu`��M��m\q�X�A"�rO�?�Ś�B�n"�E�5�?X\ ��g#w��������C�x4�
8F�^j�]G5;����Tym܎)���44J�tLxfV��w�ތ�+��H���$CS��IO�N����yږ75�,z7�HR���Q������pn��)�_񦭊���z���w�)4ſ��z�����Df�J��kW�V
����-�O_clo�/�ΥC���_Z� ��!og�3��.�g�v�:�볤[��<�(��@s <�r{��.w��=�,0d�E:!C���RO`E���G���q�$D�k�pZbB_Ğo�2�'W�P��?���9f�Zȋ�Xcf�������n��P���_
�t�%�ѴI$�K�օ~��Hº�*Tr�)U3*J���5��}i��6���R`�^
�$s��!%���<�A����0�@�${��� �E�� �D#�Τ�v�zY8�����=�	���9qY�+�m'��R�U�䯴F�o~R%ґL)��h~_K�ʹ
*zs�hUϷ�ENB}�V$8ߝ
�@�i80��Q��`S��A��#RU8�e����B=~��v��kw���k.u���c��X�M2�C`��M d*��f��2�P{�h4�sk��L�"�F1�75��V��r����Z��h�����iu��5]Mᡰ"�l0���_j��;E���l��E����r[4B���'�}����1R�B#d�?%N��������Ҹ�=��d��}W
�k�>�m$j.l	��y�;b!uI�8�U�#���(w��.u<#�g��pqN)e�Z.��r�h��TMJ��I
�WmS��p����X;9��D�aud��t��te
L��_B=S'䯝"4�@8h�	'���mg�٪g�L+b�iv�ex'�n�{���k�@�p��"Y�㪓ꪚ��J�􍈞:=zE��3~.|�;I���ښ�o9���������3d�������^��mD<� �<����oJ�+��H9ܝn��`#��ɮ����>*�r�J��R*��;��K��`�]��Y����ӟ��Z0Z����F�jM�oh�� !Y ��NTx�q4���+��c�B�|5�݀��P+A�6�ڦ7=�q�(�q�?

�LY\V�J���-u3�ñuH>��}ƥ4 ��E��4�}1� �}]�-Q:��Ӕv��l��ݝ�$�Ҋ�^wkd�Ӣ{�|E3��kcRfQ,�i!p#Mq D�hِ�-���,���i>�qHA~B�9#�0�f�)ݺc�n����b=��+�Aq�A��V��wR����o��!�T���(�=�������ғ業��[k؏����O',����
ax����L��\�B�
}μӊ��R�l'* %���3]���h����k���oV���F�k�~%}}�N�z��5�I�i�oMh��Uz���ȗ��1���|�;>n�|���'� ]�R��Z!k�{[ ���$�Wno>m�����(��V�_N]�#8�'�O�~����(8�uLDSx�u�
7���:[":
X�Z�s�qB.F�UM�����}���'�0� Ѕ�v�eVLs����	���Z�̡��LN�Y��fC�(������B��R{'�;����8�n��
��Б���i�V~8����U�-g�5e[	��R���!�d����:ں�<H(;�K-.ʂ��l��?	���p(3�]���%�n,����IJ��lKj�������'�-&!��B��A�IY���y���vL���HԫJ[��_|cإ��ARe�4�dqK�q�kt����VHK$�����_��e0s�z��F�;,�^_�厄Z���/܀z�6�H���9�/����)qR���cR���v�'�I�(u6u_�U�$Dz+���R���q��ʨ��Du�%���71e�>H�̮F�bu��jXkڤ�a$<�o;�Husb����VǙ:3�����É�KmL��e���P n��in�̷t-柏�Q�\�+��D���W���,eǎ���;�O"�w��[�@cDH��4��s9і4\+���z� �z\�5�E!L���|�-N|��SHi_��,/Wtg�ڵ��0ZjC�ȧ��ƹP��,8�8u
�^�7Pi#�C�2�blt2�|渼��C�%�������x;X��@� ���4p�?�~�S��>�ڼ'd>����w��w��PaWq�c&ޢ�A��}��g�AW��*_���Q�)�]���u��z5��v6_6�x��V�T�a/� ��M-a�g�>��)\�-��)?��O�FM{wX�:r��e��5=��I�R��2o�<p�d�@6�ox��~6/k��2��f����@DT!�T��d�q�(gq	o�v�2]����&N|�!:��VmWߑ(��XOe�xw�.�P��%89�)��FFErf��L�	,�1D�PIj|��k"�%*�Z���2����t��mb�O���)��=.��Y��o�w�������RE����d0Q���Bv/�u�ǖ����[-�v���M @3y/��@+=4~��c��&S�3�����ʾ�&�0�z�C�Ȝ,	�V��10*)���	=C��jQh?O�	NN_��D�I0�����4u���"2L�	YqNE(�S]QQ��2�+�W^O{Wwyx��r�ɂ�.�u�H�(`��r�#b��%�|K�}r����@�"�bH����o�*?
��"�ъ]l�pH/"v�ÌN~� �/�m�t:qT�5݄R�[�U����ǫ"�!�78���-���� �9-��OR��e��]�<#@�_i�$�PL�GC�x�����<��C�8K���7���ja�;���aՆ�����#�|ڢ ��b�O��F��V��і}oú�b�ۄ�4O����~�������ڛq�&ق�^�H�r���Af�G�K6네�`���d2O٢��1	�s���p��h����|L�d2��00-T�_W���S�'	ѵ�=M�K��ta��8Iw ��Oϥ����$]A�JPN���ɍտ�·
�Of?5�����w����D���a�#�����1k��y
(�M4*�ы�Ym��[�������"�}�����j�|P������ޖ2�e������H��F����B���5E���9���Pˤih�L�6��G$V��Ρ/�0Bd��ړ�P�v�{=���D���(�q����s^�a-�ț��?�Ǯԋ\݊�Z!���/r#��\��ROv%��i�&�����������DT�����)�q5�@�U�Q(�&!�]Iqp�C,����h|I��:�ٶȽg�f�F^VQ&[�	�J��KV�3-�߂�ˎZ��A����E]��0D�/gʭ�	]�UߝnNIp��D^�� �;���7y�Jg]���a�����Jm�]�3soh�yYқ���br�H�W�͵�JDe�Dfv��`�)ck��:��֯���3���u��N:�9C��))q�\i���$u��ӂl'�e�w��T�/�S��I1[X~��ݨ76m���?Z��m?H?�n�%v����P}f�F�j8����L =�lpmՒ���Y7�yNH=�T���������j���-�s����,^+b�����N��O���E��n�
`�|�*a�z�X	��A��=|`���&ey
��ʌ#�]+ �.&���������=���f*��l����g%��`{{�1��s �3��"�4�|�
g�:��PT�r�O;}���55�P!��?In�P��r!�t�8N��wN��胯����@ډ`�4����T����E�>A�F=����3ޜ�e�+�� �,�6�R�G��pL��\�4g�D���Γj��uu�S�qI�d*�P��FK���q�L�ު3��y8�ᄛ�Q�2|�h-E�����?����`~"��f��N6?s�Y��Ec`���Α �}��*�>�"��+��+���p�yq"{k��;H���[8���������g����Z�dY��
��-�_���k5�G�T����,���&O�������������=�"_��ko���@��L>(T�����Z)q����<B_|�Lc�d�2=P,(lXI $U3BD�ߞ���!e���y0Ս� �>��^)���_��:��3}���(z�<&��T�*�>n(l=�#T#��~���lj��J_Ϫt�/Fki��Q%�$z�Q������;�����8LM�b�*'w?S�����T���tV;t<�w��vf�G�vQ�}��᝵V׷p2��4�$���,챱T���'Սj���� ��1���#Զ��t��/>a;�-�Gh]�`��>LlT]/�k�h����J�d]��7xr�����/��
Z�t��o�({��dND�����6b-E���
�]����Zh��0��'3Эk�s���O�u�I�@��:a��P�A;]�R��-���M�������t�ʵOI/4$�\����gL`�%D��Tϳ|�Ke
�f������%ڪ���B���sTL��Í���&1�4.f5���X�n��O).��f�kz��fb�,����3� �(�Yܭ�ƟM�d<�5M�i<��H<�Ԟ��1�=N��6��5p6F�U�u�0�N*��.����[�2w�D�����E˟@�S]���x����p�x����;eP��3-͑!Y����S��w��l�s�Е��ּZ��������
X�	U"���f<pf����ؾ�9�	X�� Έ� n�\�~X�i�a����<3(�#���LD�j�&D�]5�SI�?	Xל�pfC�5����%I5K����;�^��k���0�"5*�-/��[@x�vs���e�{~�� ��Y�̡�N�c�����hT�H���H��B�*��S�`�L;����cEc���s�/:��=p��F�:yFrB��]!�ےvb�${�]��.�����uO}X%҅i�M�%��{�z���� �'R��&\Vԡ9��w�+R�n,����E��F�x�~�e=_���-��<���u�*��|u1���ܶ8��jU�슍���F$@�����`:O�:̓A�R#Nz՟�Û@<Ђ�,�;��ly��\��8v;�`}U��R�#]">G&~ּa��R�&��K���k����D�&������	��SH(��� h���S?��poxe>1������u0S�����/J�/)�H$.�vtLb���	,���a����<���vOw���c!����=���7���A�iA"��"�`3IY��d�P�T�ʈyk�|���鑠�( 4������������#zc��h����t�L��Ӣ�e؉*r��׺��rJ��=@a�Qtϓ��h��^����杍T!������Q��&�[^�̐��Q�p
⓫��r-���|�W@H���D4��5�`]��<&��c�b%7qCѝ�)���'񳸩��2�i����2��T�Q��c�p	�3��lߋf��d'v��qC���A��SJ+�bA��2��W���ih�!��3$�N�Id�ӵ���#��mA���[��D|0e��Vi|f9P��<���2xb���9׼�����������[׹�'o��ؓ�\}����i�Xխ�:�^Cu���.�[��#�t�0��M�f�$A�9$싥E��\�^��o���6��1+�	���\4V�!zqi��)/1��,R��^Q\��mH�!T�\Td>,C-I~��L3���mq��ܽc	������?z�_(��X�:��`%�*��>2薚Ff�ŤPlfj臤�������BN	4T"�U�1�.j���2���ꏚy|�3���-
Yo��4&Ͱr��!+�r�3ݕbJ��9��������z�������~�L����P(�Keʈ��;�7~f�9	����u>���{[T�ZϠ:�q�y
�n��wY�+�I�Eu�oBA���� ��,oj[u*���]�A�o��/�'>K?q���|���Vh��7��$Z�D�R�Ę� �k�bgL��k�9��*ӝ����^���P������ ���\�X��k��m%�tb��X�F6v�s��8�!�kG�h{l㹤�s��E	�)6�S�4�}6'�K���,U&��]w"
p����­�&��z&)���^�v��j�iX��s���3E�T�!h4�?WK�H��H��x�=.���o�qw�3�f;s�V&r9pS�8j��g��%�F����6a �.��㜚��_��I�Iv�l����U{�+~�veSߣO+glE�_�X9@�XA�]�6Q,ʒ�}v�q����KQ�^�x2N_��m�������a����h�]��n���\Q��MG�&���؋�8��`��&J��ޣ��؉DF]/�$A�8��1��LH�����	��A,GW2�Ֆ�݁����/U%�c����F��~ؐ[?�����b*7�.u`���1�4L<���|)v�����6u�Vd���C� �N�����4��J���aqu�=�������5����gK��z���,{A}��BM�����i��f�����rd���q�3Gȩ����t{89��Q�K��ro���]v[2�}�,���&�.w�|$��s�3µ��%���7��YjB�c�[��������y�(�k�
M>���<��
@ܙ���uB?XPe��U���zSnL���]3a�J,�C���^n�|4̔�m�}��ڸ5D�i�:�y��l*s�)Ow�9�9����i�jQ'X����`gfj��ݧ�G���m׹���b�)N���԰8_)'Ъj��0���<�4��SÖ��C?�XKk>��n5E�?0��#a_��*j]�]^@�a����:��z�w����j~������9�u���`�xѿN�Y��� ���WV��C�;�ے�'tO�]vz��Z'�H�'�����G�x"߫?�$:q�4�K%�~�Dh��O�\>�(��-]b�@S��>o�G�/9�e�u� [��'$+}�Y��	͞�
|��g�Z4�`���*7��0xɶUT��L`g˖�48E_h�����$����hq*f�ѣPAV��84,|�������N?5�J�c�J5�Xzia,U�T4��nj�҉����S1RT��0�p)����6SRQ�ʴ-�wh�p�?���e������ ������akn�k��I��+�Qp1�W���Vr�FκsCjBB"g�$�[@��D����3�>~����zY!U=���!�,�]Y��I�G�s���#ϣ&[F�́ �����4�Z{�Y��֛v�G��ͬh�)Y9��RJMx#�6����x�;b���X@߹�l��v,�o�aJ��dW�PGI�g�6�j�X׭��h4��|�Z�/wu� ����f���!/�qF��wN��ٵ�z�m��\O�+~l�v7A~�+�B�M>@���y�6L���o��غ�J<���&ӓzs�b�����gY:��2ȵ�'3�ٕ�� V��ͬ˵�)�����{��M}zj�~�}�&ǒ�g����[�N�,~͠�"N8�6ӁL��op�uzE���o*-u��.�jM@H���
�y|D!���W��{��'w�i�an��B���]*��\�^�
��G�����c��wۉ?�r<���j
Ƽ�����?>��O�
&Ⅻb+�V��X| �+-���kz�uIDr�X�{s tڕ%aF�"��`�~QH�� ����H�9 �[���\7�O�z�^�C+Q$Ȗ(<�R���H�@ӭ�M� �ڣ��S�o���Za@����/�u1�y�hO|�j�@�I5�tג��\�-�;�"�����')�f��g�n�:"rI+ď^
��ݕ�5�M$Y8&����t�^��=)W
zD��"�v��n>��+�x�D��+ԁf�hf�mur�s�}�z��4`�u#�0�3��������O.}�~��с�����ؼ�}��fxAn-g�^�5]u�V�`6� ��Q^`�'`z�M|���G*��1��.�=�"��pL�q�NM97�D�gzF89����j�	�:�W��R�MCI�*�Y�\��I��c��
gH��UR�<�l��&�L�j��|0� ����kop#���$���{ LY-�k��b晷�	��~��)�m�.�:b��g\��/��O{3����R��؀9>Gg���6Q�x��E�X�`��N���T���Cˢ �s/h�4)9-}L���4���궴���K'�W��>���wx��<Qh0D�$�=?�!�N^��G�d!ɗ0jK�2��k�7��pj����8�rED��7ہ3^�%�
�N�
]��!��]�Qر��!��L��5�������7Wf�plGդP����� �o��&����y0����i�ީ[,���m�0�
����@���.�'1=� �@^k̢G���-��2����h�-�R��Kly�}S�q��G�s������30�$���|�@O:S�����#	N�KY#Z����"7��E�ث�nF������D�NU䢊xuV�"��5���K�-3�(0So�)��2��OY%w[�0G��;�m��;�T@��m[i�mi���n
�ؠ�����}���eJ��h�2%^ʁ���Z:���iH"��c�cq�"|�B��2@{MK�/l#xB3�\*ﮛu'$��!f�U�|i��E��-�Gf�x(;����ŇB4�W-����m�Qíã�׎��LW�s�.����/����p�[����YL���j�խV0Q�*�,%�(1A��kgSf�����Ts��*�e7�q$�kK5��T�����s}�o;+4�R^�v�����<dI�ۀ�8���8�bk���7�0��1:S�ĩh�?o��^��Wށt���+h� u��*r�Y[y4��
�_����[��ˣ���?�w�K�*���3��\n�9]� ?T�A��v����E2笶�Á�e�A0۶h�.^�8�Y��J8�/�PA�4b?�ԁ��j|�l��~����b�\���g��>6t�-[��[\��@��N�x����n�c�%W-X&�}�a�mY	~���r�e'V�R�*�g!�v�
��7mSW��i?	�s�r�;�hl��EJ�zQ�����l��2�������s��5x��,~���<�-��eV0��N�׍��)w��U/�e�J�N�pF9������*;O��L�^��tp�x�Z������U-�n	�̅��p��`�!C�>�M�	4���́�؜��wd���Ϸ���tv�����Ų��b(��,:i�
-15s	�Jp@��i]I�k��w�oC$u��,��_wa�v���~tg��l@�ih��kr�A��fv^�t��zE�3

	3�Q=��2g4�;�*n��zm�/vv��?��r��F
ڝ5�0#)�{rN�"�>���S���H�K=*S�HN?$�*(�Ƚ"�R�
A�L��h^�r�gGV@��W�Wے�:sLI�Gv��x�WR���*�ހ>! �w&<Ć�����m�._��S�?:`�یt�W1���_��-�+~�B?��<e\J)<���ǈ�)�N��H�J:�$��e��X�)��O��}��dܢ���A�����8T�z��c�H�`R�����B��B�z����s>��`�W�A��X���̇�Tv{���w�q8`���ǌ8�����)[�]��#���~b&�x��4����a��.2Qvi%e1��q>��^�,�FPu�;d��Wy0 p¥��R܊��B��u 9azX�0r|�OW�&�`��_{g+���X)�ם�X؀���a�sP5[ ��g������[5W��䘆�;��c+{!�K
�wc�{d|,�-y�%�7�ط� ��9m]���I�{�&�<N܆j�M\��@���"1�W]�g��Βw�s��R��"�d*�
�$qu����VNۄ���[Xf�N���|<����{~��m�������'�� ��2К����oFyd�J�`W�ab���tU�'��Yp�Y�4c�7���r�ܚl �-�Pz�{����
�OO��n��AV���(��XF�nW���TE"D9�<d�!V��:��n����I�$ޤ,e��{��;j�v~ߩ��|��8��l:���&ў����'2Y��7�n�)�w���1:�,R�۰���n�dgի�wy�('T���z(��s���5����W��RC֎윞�e��C�p�.���|�6o�\�b	´�Zq@���o�G�lr�%s��@ $�%��#!
,�$���1�Y	IFl�|��17���X(ve2YH�HDv�$3=����4r���jN��%(���D�9�ڭ#Cn`�c�����6J���PD�&�^�fA�=f�{�����/�k�4J�,K;��Z��>&�]Ca�=É/���G̗���^!<�)aMC^��}����u8���!�a���J����P4�q��LC"��g3>'�I1���է�G�s'��C�@��v|w	; ��o�ٳ�ӏP%(H|Sef�A���RO{<�}����=�$��ק[j���1���@��g��T��sO���'w�:Y��z)��(~�Z��A�1%�u��B��������6t�p��n��3#���{���N����f�/Z,`�(�$@6���oo������nk�5TsP����A[�|m,��B�]Aa��������3h��� /ȩz��ڹsrF|��ee!56χel�>�I��1�;���@Ȃ�����H<�KV��|98eM���[H��Ë��м/�>n���bg�+\�I��'�3�csӚ��� �/��eO�d��99�1w�]B]nF&4B)]%dd�7/>@uG-JC���8S@4s]��i�$�3mt	$��Fb��`��:�0-������&��4�He�Y��Q?o?a�@��0�0����i�=49��4-��n��_:���ł�v�����Gg��!��c9?E��p��FZJ�W.1�,��6kÆ��}�J�!�yom܁����#�?^�I�YV|��A�6���3�(��$����� ��2Yw2��_��I��Nzp�t�ӓ��HNۂ^D��;Q��	�ƞf[˃���Cx�|jt&�u��IE	�C�	�5�Q|٫���3���s/r�E���@ �������f��&��3Wyu4�#]H�oi".�ƈ11��،W���u��7賩��Voh2�?z�6�[�|?pX*�VC<ؘ���U5w���Oѐy��N�	������#d�[p��;�*Xϼ�+�����*��?�����;�O���37^z��{�f6�)#�2q>�(�T9$Wh�#�U�f��al�;�!�A�h#3���� �+��9��6�PCY�-{.?����<6O�5�+~��R$�eN~M�J�l�xB�F�g퍬�^����Z���7zL���Lh1���"�0<X�3(ن�^�F� Dg�/ a������4Cl���*�\�����/��(�=`^�Dq���W���&/�𚺆t��w<�r �}*&@�}(�����t�Bw^�i-d��b��K~}�؉M���ه�Fn����'���ab%F�0�^|>��ojsj��;�0,�3�#c��E�vE@r*�a�u :����4\~�;�93p)~����D����TVޟ/���2��䢾��L��T~I��Su~�7Ք�
�ڙ���m��嗺$��3n<�d��9����X��:.c�᫦���2[�^���I��(��[
i�����SUgC��+��]��7���#��D-�BR��l!�$S��Ō�[���=�j!Z��"]¦��O�������󒼭{<��=s)>�o�3��/o1w�Z_釞����HS[/�qڻH	BR�d�W��~�U' ]rW1Y%��4wrﳶ��y��8���w�U ��Y��Ǆv�o9
�m�A�r���_��o��8ށa&�$1j\�q����r}E�?:gr�~�4E�8�:^�(�'��o� WZ�B�RF�Yf8�'̄^�F!�@�i]��+�>e���=OWP�<;:�Iq冚]Z���!('�/�t����*}vi ԽaF�bA���rH�
pkdڴ2���� Z��=_���UA{����(�ߦ���#�����<��=v�n��kh7��Ȯ���L��+!���=�d
�u@� ӔZc9��@1 ���.�Þ+bs5Z���^F�>b1#� �\�ro3��҇L���u�WK�Vl��:To#3v-�o�d,��"6�y��nA�������A����@j#l��+���2��{����L,'��ɨ+C��݀Rz~���U�i)z,�ݫ
�l���_������c��
�S��kp�M6KE�
c&؃��J.�I>�6x��n��@${*$��g&�=�>���B� �<i��Ń��^���=�MJ1C�yq�H�^�O�E����Vzuܚ��������Hx�D���w@;l��S���g'd�?�?��E���SQ@��\�p!"'랞������ʠqR̞��i<�椦6��E� �o=�I�^�I?\����p֜ޑ�i����1� 6]���^�hw�� ��c�dtj�)q�������?��%��H��8�{Sɍ`V��;���,-M��~@D��B��7�A�����)WB��۞U��FroA�9��ͣ��U���m�8/�&S<�\���X�|��=I�!�PʱS{F�H3�Ju���m���UK�6����FԷ�.�MI��'0�n%X�!b��1����"�6t��R�a_!�NؖX���\���B	{qƁ�3g(YG�tX~��{sbfG��+o����S�mv���x����+d�M�JG?����ȋ�He��ep�0�KޜM7��5=.�L�F�eG�������άe��jm��d��%���OoJ�~�je��2���&a^$R�,*���&O�Q(�\y����!M��V�eP���<V�U�!�Tm�x�t/�q����H�b�'6@D�_D�~F��@/`��0�;o(Ȍ�7�Փ^������H��-�r�/� ��ײ��<F�I��lv/�
���ջi��1[��zRU���.�����4��@�����
B� �-[�����N�~�4^��W �
����K��z�LX�0[�-I�R��p��v�~�"��l��P�ه��ih��L��i�8����]���6�1����\��Êkx���_�FZ�bhZHY	��[�D�W)��]gHϠ�n`b�]wSB>�����x)����O
��$*������bv*uAKۈW���/:F+�QX���oUX�a
��Ԗ_HcGd�v�Au~">��&5~S��K��1+�Vn+���R8<É��S�I��،������)l���&F�?�GrC[�П� �M:5b�K� ��{��նC!��^��\��D�r��]�l���	~�<3��A���|.��b\�o�Wh7��S"���߃���u��f$@PUꮸ��rv 
�rZ���w�XD#@8�z�6������v���B#�O��̕�R_&\����"��+2%�UTb�� 떁5�3۶JΚ<��BLJOu;�9��*�d����/�<\ ++�}��
*E�D��ٔ-C�p���j�l$�=ӈ�� ���B{��؏�C
�ͱ�U4{�z�і�u��s%$���1�]9��n�s#��դ_�1׉�h�����=��H�C�F�/�.��%J��T ���[�X[�eV�b�l|�)���2��7"4�j��ݩ�z&�$���������ZtΣ�ZҌ¡\M��(q����'�ڼ�zXQq�O�W8�p�n5��§�|�*��&)��ɮH:��{���aב-��}��W��W40�9ei�
o��|u3'�:]�B�4g�AE�� WBe�mx��;�mj�����r�ԑ����8=1lH��r�i�[���p�N!�W߿��(�7�1C8y *9��� ñr6R�| �6�EU�N�LU���ETQ�̝X�v.��bc�U�,�^������a�>�4������7��/Y�"����T�=	Ph�~:�љ7`�^�K�r�#��fp�D�h�&�R�WL�cyV�T��ܝ�u7�aEp)�]j�N&wW ��������KT�h�+������g�Ԕbǘ,�����}jh�y�_A ����������
�Y���
�����5�;��5��&�z��q��1�47���r7�gv�����\�Z�Mr;pd�2K���I��GO��xd:�At<0�F]�{pg$�Uj]M����s����"{D�[�%�	9Һ�u���H�����Β��CY�MJ���ԅ�bJ$T���-hR���������O���4s�^�B�J�k���$��~��_�|�^���R��h��S�&E��)�HƑ�_<w�j�L��H��ڝ!�HP�&��m8R���A_�i����J�����lt�_�ԼR����<��s���7���Ɵ45E���m��O	y��*�/�t���`��~�T�[h��W2�0��N���ҏ�y��q���%��V-9s����I�5!��<��J�2kZF��ZJ��C�B�ˇ*:�Y9�a^��dS��I�
.1vѧ�|�w���	���r��D(�s,v#8����K�<�� ˇb�Xz\��S��`�d�x��&����x��>�1��3���^��\S)���??{�"���Y��y�J�~�i��U� ��x�)9}�\�F4u�F��H��2�	�����:�GL+kG�L%�j!qG�#?h���V6+3�G�ۀfe9�No�H5|�^�)<5��[��;W��蕭z�U|��%���c��\u�������N�jڕ��*"��,�h+T6V-ɧz����i�C��1!�����F�4�Q�.�e%��2�7�q���)����+],m3��N�h��/ܗ��spD�zz��y���H!9g>b����p�I�]� w#���v��P���obz�{������>�@f�X���W��Dv�O�Z�K�$з-��x�vԕej�y�m���g<`1I���'0���8��� A�|s����� ������M���8/�$�N����)B6	��W)�D��Y;�_j!��{}t��h��K�������џ�GI꿐�6���a�K�����sH&��+��]x�¡�Wbc� ��G����l��xO���׵�Oܥ���B�~y0��?��C�u��2�М�5�%�Pb�a�/�ܑ��THX`����諛*eT��@��ҙ�0�h���c�2�x� ��礚A�E�m4���&��'�M�v¼��,���8B��t�7�����}�������D���!�����T;	WˎOγ9�/���!���:0�����7�%����ߑ����J/W�ŕG���_���E��BٙP��o��EԳqí3�!{n�ko�&,]��$�����,�Ր��%�B �M�,l�@���,"P|v�g��u�?8"�j�7�0�M+��-�7s�$������}���3-�����|����Q�p���[����f���g�3#�*eG����r�-�T��	6i�B\�����*	�n�&T�D��/+k&�G>"-�j`(���c��}�7�0i	��ޅ\��Kr���Kh�{�6k3�����-��W EW����u�)���/�kd|��&f_Ţj�z�cw)zj.���0���k���<�ʊ��]=<;��T�hcb�X���)� �{�����,ǎ������A���z&�K�� �m&BH	�:Sv^����fv��&���E"�LfD���s[o]�f�{j&�z��{-@)�#}�P
v���o�ن�-�ë�(�����4)o��^^(�W�)�R���V{�2o���]�D����`[��#�*"�˩�wb���↚��-�K�_O%�؅}�<u� [�8^L���ψr�2�ltJ�.��I�s�Q�f���8��G�J�Gf��}[k��ʀi�[�k��qWt�/`�������:�O5)��|=x6�4S�[�� ���z��X*pV5'9���3�B�WE[k�wfh���1ق�H�hmB���3̳����n찇|GE�N����c>��#�)�O�h&�m��_�1q�e�-��
��%^/QE��܎/��GgƷ�܉��ťb�����E�N(��:Y`-\� �v�y�1�n0�0�Vv�+x�B;<���7�����ոߩ�	}�^֡ўIi�?�݈w�۷I�#�Ұw[��Ȃ��>$��L�@���ذ�
���D�?JN�v�ER�mm�	eJ���g>���6b�c�Œ[k���q��I�4�S�����W��!������?2{��W�K�X��I�QO��s&�?F�n��Y⨟�/d$��S�"��5�8~����-6Ⱦ�_'���Џ�/CM{����);+��]���R .Sŕ��K¤/5�XI�����k(�
��jn�����v.kY$C��癉�^�� �ڠ�~�����4?_/юdu��މ3c]g]W(K��]�����(Ԗo$%�{����=��x%YK
��]e�D�V]��e�ђ���r�N������#3boH�p��[�7�8V�Hpی�}�х:+��noҀ� �k���!�8�K��"���cm}<Kb[���]��y�)�\|�]
~�!rm��ð��V�/��=v�O%ʃ�U�G��ۊ� ��b���eZ�1��DFOc

 k�긅���Sd��X�r��!���Qu�t�ܜ�Ր�8"1H8�r9��LP0 .^H��H3�(�B������5	�}ny4Y7�ϖ;����ZQR�F�K<U�`t�g��G��ؠ��ӳ�{o�R��?�+R:$�f�����,H��Cl�GqK��>M�)U3`P��&d�xf���?>�[H�s��n^�؃�B~7c$��F���+�`g�id�<�]؜�	FfzFLʓ�b-N��a�:�~�x���2a������������U��m*X�p~8�����(�b����5��Er4���N�>�
��32冇��3�`���勴O�٣�q�����Oa�������B�5t�ƵN�ZۦA�}O����F5@��e�iYb`��l[���LQ�[���&�X!��H2�׼z�k�IbKC�4'f�S��ù�A��{�N ���q]p��F���P�z�'ԫh��4��c���e�x�(�d�6���ӓXdb�#��֝Y�m}������`ع��>��Vv��껡$�E�n��7�i��$�{^�G�h�:)���]�P�(X���5i���P9�L#�W:�M���Jۆ'��1�PSp��	�D����AvU~	ۘ�"WЁ���r䜣D�Zc7޿Pnbo�`hJ���lǈB�`��Bhz��B�<���u%�:Yoc�9��WÚ�5�d�B�$IH����npV,�l���T�D3k�s����m�Qc)�Uʎ`x�� }�R�T�B�L��&���%�R���/�8�⳴�x���΁]b��k�](
iRlo��I\W��Hۏ�ꂂwş�j��-P�T���tRX�!�3�PRJ�-6��4�����Bp[��'B\H�;������h� 2]�zΣK|�\��'b��%�{�ކ�@o$�ӑ�;��j�`QT���tfT@��Pci�������tA�뵮Wv`��?f�#e�˹��{p��9`eB;H �W�6�P�����@�u�rU��9,�0jTa8I�WCӔ�ʻx�tmP	�Ԧ�E�$�5��QK��Z�R ��&���/E�՛�'��fC����9%B`��pO��jO�gdv��{�CW_M'7⢋��M�B0~:ֲ;p�����DV0`>����T���%�gLi����fe�&�a��'�I�	A:VO.�%�+��Ok�+a�.�E��.
��e�S-!v��5bh�~z�샐�)�a���Ŏx�մ(�1}L?�{����0=K�dB�؅D��޸��:K3U|UzCd: �^g�7�^NQ��[�JX7Z�ZzQ����qv��o�͇T��P1+�EF��\�4j�k�� �0�����y���,v�JE��@WaI^G�X�3F����i�k�)�.��-�X��-�>�1�����[��D]���@���bx	�m�G>�}�UJ9S�}�s���߀�:��$��ѓN r�h�����dj��������f�9�������/� ��h_](��;�\�6���}���c'y��G��7����2hވ�n�����(��<zY���y�{��+DF�ֲ��a����_)%�p��߮)B�x]�m�F�#E��J�R�o��	��+��Å=t�R��-������&3Q��� ~����D���ϣ��w�rT	JOtuH�ѩD3�pO��T���튤�*�M@;7�-?��_��j�Q�C���.��gpaCɃuVQ�:�Q�N���R��l ԘO���p�ɠi�����J��3a[4���97R�_�[�˰�i1��z�j�Fz��J��,%~�t���4�q>T���2شV$�H�^�E(�r
�_�(Ｆ���0I�n��#���I��3���2N�R(LF�t��9G��,%A��n�:�'�d���=�����7�*���H�q+�ی�?���,�%���]o2z)���Mm5��)����p*}��	��-}�w��Q��+Lf �{������&�v���˵�Q�ͲI}L�>>�7����7�sv�{A�Lǔ���-���[����ұ.9��G�=zN��k�t��װ��Ą����MԏFZR��:�]���������oG>Jݐ�Y�AS�6�M�?_w1��e
&9���{�t����D�Sa~ "�1 ���+�-o��p��b:���ߑ��q���^�f,,/i��jUe�;"�D�������O�f�C���JC['�6���}鳄Te�)����2�,+��� ����G���-I�T�"� ^ȿ��b�0�T���	���S�������6�V)�У�w����d�PsC���j']0i
�1#�,f��y���C�fqd�BG@��+b�;PR�ЎC��LbĒ� ��XH�8h��PyF���+Q�ȟ�Iٞ����}�T�N�G"f��P���.���$�B�>t�XK��1��[�	�&g'��*Nw)i��&;��bW����� %,P�ТG�����k���#\���W�-Z��!�{D{�o2��u�A�\��c����͎dl��>��.�*U�Ο�~����,&"gJ3F��#�pIM
)�:�l"�.�1�y[U��b�s~����7��Wج@��E���0���H��ޞ���h��� �1�[�N�����q�Ŕ����cj�	K%�#��P9�
���[�I�@��Qf������Y�4H�ߪs�����5��^7�������rV�u��+�K<���_��"C�W���_B�6�Ǣ}�dY�Pq~��"��X��;�C�\y������H� ��g�M�����m	�@�U�*��|�yW�90��E]��)^�[T�򅅒e�5����o{�`��&Q-F�,?z���7!�ALӜ_�C����&;ƺ�2�A�md�L䔗!hY�3�ż���9��n8��y��"v�{?��sE��|�r�����5�DS;�ߏ�0�����1˔��۠�SѲ�5(���#g}�uf=]/L����/�����_rG&�"U���_�%��������n�p�5�F{���S"N���_Z�Pu�e�M����Z�g�˸>z�e!)߫�6	�du��l�.�-�H�����>��i�LƗ�
^��9���|W%��^8�nd�To���^e��p���\m�}׽~oөW�dt�T��1Pa�'�y�,1	l[�.'��l��>`�����U�*L{1��NO8�ݸ��w�u4\����Oo���,�c���(�>k���֎�AP��2�P�H�%������A��n��L�׮� ,L�1C�qH��.��_ ��k�Y s�/�[�w��o8q��̍�ꞳU��rB<��]���y�8l�LYL:�|�ߓ���_�ҭ�hT9t�I�l@屶I6E���j{w`�F*��@4�}o�ȷ���%b���:���"C	����,��_���dE�:��-X����D�]m<��J��d��
���Y�^j����F{�+b�1�z���H���ʔ�Jɜ�������iv�>/q��2������X2���+[�X-\.f�C-ގ��bL6�c�c.b���q\��V�t�ӣX�e�C��[�U&l8ła�3Kс�8Hņ��ZM�Eh����X�:��Z�8�|�M��Z>��f��\լ�����-���n�<
�F���L�u�I��1M޶���Զ�w�vș�}��O���s��nk�t���3�f�sO�����]Űu{d����ݾ�&� ����p����QI$��p�kX��~\}��Y�V֘�{V.\�5o�9b�#v]�c���<W��Bp ����ڡT@���Q0v3�:ٵ!	ȝ�w��K��N-�Q8��S����B��QWYAd��q�B���$_�f9D��&?��$J~n��NED���m2��֧���ˁ�W���H5����ASIB�~�ؖ�����r �����2��q��eD�{�Cx޸2vB����\��ͯ��[;���Y���_o�1+J<�G#B�b�Po�E�6�-��dHөA�.��]���I�Wϼ+NbO����d���ӊc�=h���nG�7?��Lj/k�됝���w	��jj�Ქj{|~/E1V�����g��y@�L�ֵ0smvs���u p��[޴�c��y�1�[��tDG�vb�<��(S'�?��o�^ۇ�tNl�Z*;�h�����0����{���ۃ� ��ئI�5!��p�x\6�z���K#�%�E�Е�ު�����d�IT4�t�D:\�~�� �a��E !�K��	��Uԡ���f��9�B�"h�!�BV~�U�:�v���wd\����dS�,������^���K:� w����9���Ǜ�Rb�b|�N]hِ�ۭ�Ga��Y�'J��6j�s�
��t|�LV��.�9O'7?:�+���Rۊ��m01(�?r��P��R-`U�o�i���&�e7���K�>�Q:���#l�/�6��t��|iI���<ӓO~�	̅�ˏ��W_vP��A%_hkj�����e�Hk���O��u�P19������@~#S��lU\�΢�>�Xt�I\`��U��4�;V�m�Fҳ�NA���Y���D;_���/���d�4��ri.GR�5ko��05��z���0 H�Ee�%��k"����]8�!�^ApAL8��?��*���߶��S6��5�VpI�.R��g�_2�`�[�j�c��2w����d�x���R̠�]"ˠV��7��kn��<fd����f��I�j����Bo�;Q9���%�aCN�7����Ca/%H��ɿ����+a�m���Y�@ݗ�8}�3��]>>g�0$�xJ���W!8��95҄3HA)�����|��ܠ�fR����
��,�h��kF!�ӧx�R�$5�eԫGl���=����O�}�~"�9�Z�h�Ֆޫ���yr�6�DE=污5��V�fa�7/3$������Q��K���vy*j�$�Pb���X�a}$�����Z�`:)z�Bͥ֠��^˜ϣ¶]�ҡ����z��ڀ�a5����W�-�7�ͺT�� z6''H#21�Y�;.ˠ��������@M�V�޽�/�z>ca>�SKJ�{^�4Y�<�P��t����pK�Ec���w)l(��x7�!�B��j��du�b-�n9m��౛Ϳ+�׽f�"{��.����Mr'��5ڌ�o�	?�k�U}��S�!�mQ;y��]�p�����iA}	��uA;���+�^�0أ� �9��Fm;���BIa+�'� ��-�.�Ђ7E%�5���g^������EQC��?ݧL�~C�=ա���O��؆s`�xX ��~����!�iğCM���8�`�AjI�9���Hw\U�X��n5��ܠk�ar��ʢ������<�@���ȷ�6�޹c.�%yf�*�'����4O�9���+!��ՂN~��U`p��2^�A� �+^��U][��N�	 :��J[�P[Sf��t��	d�"o+EJ�PO~-*}�#	���JŖ��G���o�6� ���P=��t9oG����>l�r���&�����{鞜 �H�| �0V[�6���U�竜���~���g<��Ǜ�ז���&�!!�g A���8��Gt�KWXZ��lg������*s�~��u�R����񢨼[J���W��V۽_X��>b�w��������oA��*!͸�:��������v��DƕA���풘	$�hP�ys��jN_�NEz�h�F%2����d^��(�-C�
}�'���)�*z�b8>���u���[l��А��a��$!�o��M�W���'hFiJT+�5��x_��:�n�
�GwF�y�t"ڗ�_u	q���� Q�s�ಇ�1ٸ��j�1XBO5�0�������>�v�/���G�4�B�$u��Z,]��4������͉�oM�Q����t�c}!�:���L�)n�=�K�I-��ȩ�V�*���ueб�C�������P�#\�d6��D!R$_ގ]"���d������#k5-Ȉ_���$�W��"�Bojw��Tw@��y���������	Y��ɮ.X����6�I!?�{qn%��ӐKn�',��j�˹.�� �����Ldx��rl�:��H�-s���0/u7������ּ$���ҵ�{N��+V�H5�2��ߞw��͞����r�sƵsX�������l����:�hT�oa%=�,�Z&t�o
U4�6.*�TNM�-��&�}��4��*y�Z�x��Y��-}؃�<��@��C���.݂�{�:2v�Z���d-�9�y]=�K|���7���qVS�Z1��{jj��4顂�G��'������B(�'��<��\bm�)���-�E�%1_�&�u�r���O#~�BA�H�9��KQ�5��T��lp�"���v(t�:��Q޻��S��Ԉ�g&z������=}8ƽr27  ڂ'nF�.�����H-�H����$�BFSd��)\�����XZ�&Tֹ4]� F���V�X*���-��*6O��ζ�/�@n���a���
���xT�pR}�&KXJ��@�]�ٶ6���yG�>L��#�&q1����0DO� ��Y���6+ZH�ϵo6�FP��� ��,w�7:-�Q�D��T�T�mF7!~lp�!��2�y���ʈuaҋx_��:A�^]@�hY�[	���yv��&��N�fAE�e�z�D-A��x�%y\͆yD.�����������vf�}�,����/W��n��K����#��	�H
�m>���qWǹ3�Œm���i�B��f@��Ҏ},K�؄�~�i�x/T^�gm�O� �v�3/��'E�Y�0�mS� ��t״�N��̣D�P����r�3W5a���D�;���@�W30��3 o���'���1�N�>�Rfb�2��k�ֶ�	��tO��o����Tc����Y�ׂ�l��|S�[�T3�Eʅ��/#6ב��.�(��]8���� ����S�ԏ�gA*��/�tk���k�8�5B4���%r���݇�)�u��ARik�*�~��r(h��;�9��ET��]��� ljHv;���ɖW<FJj'�힩uy(|j�q;���E�mˉ��6)�2�wHvqNx =�R���ԭ	7�ģ��8�����{ $������^�pcqq������j2��T��kw�'�\������/��A�3t똗���Q\b��'�Y�sb{��2'�0XXɊ��7�	bu4�X�\s��B��R�U�@�-L��0G��"[��t��7���A4U\�p)>}��p�?t�t]J���|�x&-���C�N~(�q01!�='���(�+>Ƽ.�-=�Yv[�O=5K�ː��exZ��i~�!��@�	+�XH�'yB���
�&�D&FD����uw�[�ңL8Q��cPو�5*��-#%Y0E��Zt�)e�D'�>O�,jI(�ڙ��V��m���Ʋ��0��.:�l��"G��
M�E��T�G9ܛ���:��@� "�0V��b��X���;]:=���j$���4!e`�L�x�E����#�|6^
v�[$�2~�i�+?\�n5��M.U,ީS*�j����ɍw� ���A�?�g=��+KC��V�_'���t�i�V��,[BqRS�"�.�Ӵ���8�&��ߎG�0 kwid���F7A-�#�\�{ZP�W��/%��'�O����!��H]pr4x����̊�jߚ�}���	��헙�3��.��=�gV-d���H�)ǝ��V�= ry��yd>��4�ͧ�?dbm�#��e���F�2��������$�x�S�qj����)#�ʒ�yӌ����~?[­
w1%�g��_�q_����v���(h���,�h���%�]�]*����^�ˬN5mϟ�А��h��.��G<�S��G)��0����9��l���k����Z��4�_�Q���JI�˴O-J�^ Rse<?J��P�,�5�=�z���S]G{]lҌ\~=�<V[�w����pf�z�A��"�l�)��p��z�mC�ℒ���Ϧ�l;��&{r��w2�����zk���//��)��Lj!6���)K��(��>7��֏����H�?���$N�:�$�ɇ��2r\�|�]gD�ߔJ����W*�}~YD�:���\,L�}�ݢ�����>N��wm�T���%���e7kE���X��P���S� %eX�k��[�U��#N�6���x��J�턡���˘!�v�Q�u�Xh�zuD�1�/�蟺Ǐ.����0��9|,C�6������өv޲���.�8}�&�m�&4�B���pH���rT>�6~�] ���d�`i� B�?u߱��s��������-u�� W}|�/�Ej"	�O��U�o��!�z���L�Z (�[����A����"���{�Q��'p�"0y����3�*/�	
ɽ�]Ȼ�Z7T�Zi�,��88is���ޕ?��>��M�=+���R[��#�C�y���w���N�6l;&쟸�����h�����0��ҴjG�k����{|�:A�#��W��H1u��ٙ]8�l;50���#$N��1��8d1pW�&����!�^�-���γs��	�>��ߝ(�ݲR�٘�֛������O;,4y8�k拽r����S���K˰��A���!s:=�� n }����جDS�R�@��eK/{BoN�{h\���GO�Y������O�z{�1�"���u{�O�5#64E{5?`�f��b�%���N��c���Mȷ;h�;M�����#k�P@�@.ݹ�)͞r�ח�D����'T`Z�0�c���j���5;ҨfK�<�I_'��t�4������o���?�0|Y�s�A���I�T��u��z��h�Xw�m.���]�yzw��E?<�W��bnu"��H��}�9���4����q��!N𰶈��Rf�Z���Dލ��^"�I��I�Z͘����䇯���o^a���Ƌ=˻�G�E���T�/��X'̉
3'�"z3��@)���ʹ�t�B�&���J��0V���h�@ �Sz��#i��9��֥ ��z�����ѥd�G�*M�y�$��͟o��/h�:i��DեW(퀏$�㇊`�u�t���Ȗ��銑w��4��H
��HΨ3|wr���2`�����K�QRuo�%8t�ԫ�0��'b�.��ؓQ2���{�>y�,+��	�>��R懜\E�H���7�_�k�C6�e$7��2ڡ��!�����	MZ*X��~��{��),�P'�F���Ԧ*�ρ\9/��}/��S�PXEv�`�+9����SVaCL�V�U/'}���Qd�M@���en���ķ�� ��C��9��S����B�M�5�9S1���^����L���Kj�mA���u�����5eg�,�A-���/�~$�xj��}���&�x�s��v�nP=6��L6�K�O�eZk�qs�>���"�Qx������HC{"�ӷ�]��E�����F0�*}�>����!�ￅ���5 �f��C���H��C�����h�b���"aY�gD��)�)�mU�z�I<e���!��IH��%u7Dw��2���]��Xj噟�a�*�R#���g=������V<R��s�K�كo>4|�zI�c��B��v�0�~�7�����Y���T`�U^h���G�?um"�R��Z�7�/�a�����z�����(ߋ*�k~��w._����B��ᘳ�d��S��>��C��'�)���j͐Kü$�L��t���$�/�LN&?�*��^��b �d+�m��&i뒫�4�B��R��ߋoy�ԩ������X����T�f�>y�l"���k8���"�t"�/O|$9��ο�g�3bU���_�~:?	�\9�B��Il�.a�R٫��}��KD�6���ǺW݊W�>x'k��FtG�+�q��l�Rd=A�;�2�d�	�y懌�v����M��.zj��`i<���o�R����"��o�k�3
}�b��������G��'��5�ǿȟ�USX��q��?j���l�WS�٬� �����O��/���SI�Dh)�o�z�)�3�:������/��ե�r����{Q	+P^1�P�tO1���{�%�;��UcKR�PY-bd=i
��҂+���� �푋��'M�$-C-��CҤz�q�2�J�P�Hj�ņ&��]6S �nAհ��&_��^@��v@u��3�1��Gg�K`�X.�L̻�m�5��}6�g	I�$��+�sz.��b�����?����1�R|tDƃ9X!��۪��X�S �j�o��S='�Ơ˧P�v[W���&q3�i����%=��@*v��	}� Y����V	�t�����L$$LF��=�l�%Ѳ�jA%6���!�J:��'}�T�>�@����ڱ���@��9�sA������7��8����C+P���k�WTm��^.3���^�5"v����t��\d�0`�b�D5��'	׺l���E.Tg�;H�:�v�f�P��ǋ��/pD;��S"gi�HkA'�Q�o�k)@��������8'UVC�� jS|e�Z��ۋ(��j:�8�j"�7����p:�|u!��M�q'X�lȰpN8CPx+FBis�����Սp�B�����1��<Gg���^��$g59"r(%n�)�┍�^DB��YlR��oq��ӽ�/A ]sG���U�,��N��*�B�I,B3r�u�-<�/�o��NMW�l��G��A�^�6@w��+odͩU���V�U���iM��\��^�e7�?�����d���$���=�������IP�H��#mg&�W��`"'mo�-�^"����0��!��ƻ�3A�@5?r�-��s����݅U�&Bp��M��/;�vx)O1^)~�u�k@�DH� �d��y�3�>(�l��p$���k�����1	Pq�;e��3Ϧݨ�|.���>����#���@{��Z�~TY��[���y:N�Vt��yFd�}}�r��v?2͵�����>�}��&���y
Z2:�<3���Ԗ���F�˫?�Я+X:-UQo���CMU�P��eL<�O�����S�+�C���&�l�?��"�W�F fQ|�i�X�s�F_+1��k��3M�s�mn.^1�g{��H%q���h��7�S�Yj8BQm�ņ��'v������p=�H��1۰|Mq�v�x�8X H���;�
����E��ɜ11�c����򚦀/[��:�[q�cVu'�r?]��bd#x^�Ҭ$�԰yb�-�ɯd���b�,_B�[���ۡ�sKn�5H��B��������ſ����#UfJ�_�ח���
����ÙAp�����6J"uzv�n�k\�g��L�PGa�N� t�ݔv��sc8��	7Ƅ]<I�x�y�����ΎYӚŕ��I;G�>6�?AV]lKd�������H;��� �_��Ǩ)�r�?��>�)�`�H�%�A�&il�s�Xa4%�(�`�e�����V�d�f2�Sj�����BJ˯~�YҾ�Uј;.<�	�b\�0��̃<�돔��9����)g딨*=z��x�\������93�_�Y�AQ�Xǈ���K<p�ׄ MU4Fո���J�da0:�´�l�@o{k��������o��n&�����p����o�0:G�,J�K,q����#�z��-h��&�n��7���u��bM	Rך]��@UlQ�]Z��Z#�z�w�H�L�)�=�W*R��W���2��䢶/�CK�wÎ���T�Xj�y��3�*��
����f�B�Gj3	�A�qW�J��b׏ܗ\;��j�Brd����VYҜBI�B��J��.Ҡ}վ�jI���`��o">��R>�Nh�ؼ�Ԇ���bi�:����}����Ҽr�	T-n���$��k�(�㤅��� �_�l����1<6������.�Ai��]@D��U��g x/���^��rcjn�7F�=�t���s���#se@���Gr��uhRc/�1IB���5U���m����>К��h�͜���`����;�&������cp9�+��CO������N�,m�0u�Ъ"�@��D~�� �~8��x=}b*A�ogn�����^��������陋�+�C�������kzI�_���Ȉ)7.�]y�{���T�8�ެ�]�u���y�)�������1(�1��/dZV�����v����w��ͮZ�?���÷�,�'�k�$�T��9�on�e�U� D��K�.��($8�ճ�.�=�ï4-?}�̑T��Z�P1�\�#kvѤ�,�U��U�
����"�v���x�1z4Y�oo�P���������Y	�BD����*���%��g���/���h	BW�����MHO���T4�1	�;^]S��;hۂ�{[a��B��^�6Mt�_��O�+$h	NI}��p�D�G:�R2H�E��R[��ef��Ԅ�
�+H�C�V��:�{��j뤼�ưF���ި	6����eҳ�e��[�P�������Ǝ���^��}q%Y2�t%�$�a� e�}!d����v������-b\��I�_�?W�@���4�E��M�H���@ed�p�G.J|�ݖ)��3b�L��[�Fm���A�'�hl��GXC�7/�lz��C�7i:1���3O���{��Ε�*(�������ܽ��/W�1=^L"�F`�nu���Oz�T��]/�9�kOtC^E(��s�$��E��J�z�������S���Q�幸�`��ȉB�E��Wx����!YD��b�"z�w�EIvx�Щ8���!��כ�5�C���f?�0
Rqu��J�+ȿHrUv��zB�K��'������~¨䶦�4��,h髾��`	 &5�_r��x}4�)�K�SP^��^}�,��Zy�9��o~���a{��UB���V��Y�RJ/n7�q�T9�ƨ.j�3�E�wpE�$6��t1�K;��w��9�)�j0�č̮�{�@~���A�i����kS�u<��a9΄�he��26^��E
�c��� A6q��Z3�p���U���R�@�K�;؍K��K<�>��FI��U���bE�	*-�l�������CHLB>�H�c�)nB1�ʈR	-���N{�N'�_�����"�w�	tcf�(cΟ����WK&�t���R)R�mK�Ԡ�Ξ�lus��Q4V�۞jz�e������`|��	bx�~�O�H�;��dL�rj���.c��w�i��Y��ASk-���������?��yF��%}A����Ʊ�	���N��.}*d�m�/V���x�#Yt,$5��&��=��Wך���Lݏ��Au|���7E�j�D���Ƌy�����c�0N:f����0�?�T���gf�����D�Ѳ1���aRo��K��1���5�{�S�7T���Z81�P�ġ6@�U�gk��=ˊ-�^�̹�l(�+���x�n2~��ϥ�7,�[�L���RQ��Te��zj��ܖ^�����3g��.��9fX��.
�Ө��m2��QPW�s���%����)N߸V��Z�����g����u�p �u4; m�vYL��� d����ݗf2P}t�z��	X
��v����!�A�����|)�㝗�F���s�3+�e f��<\*�b1d�Y��eU�tp�����_�~�{�j��<��w�g�C���S�w^���T��|��G�F����¤-�zH��R&��#*i����\Uc~�x�- u�u�%��6�H34�o�geǌ�3��S��&4U bq[�d��kY���}�Z`�C7�O�@=����{�t�H[	��@���08��{�K!�ѱ���A�xY�l�@&W9,��+x7���GC=�yu�h���%�u�jV�&|s�Z�1�l�[��ˢ<�|z���L
/�s�O�h@B:'�U���o���`,�n����G+�����s;�G���&�x[ƙ���X�5���-_�S��-�3�e���|����R�E��X�DUE�\�s�m�v06�{Y7����FA�DU���~�D���<�U��n��,���Zb��eCwݮ�l
v�$��E
pm2{P�L��p��5��R_�f��$Uh�^���:���=�~D!�)���_�����f�о����QC+U_�^%�B�O�ҹ��hťqE�;A��K>�m��a�3xdev�&2��d����m��'Z=|l=霌=�"P'F�\/�0��j����pO���x
�E;�����GE�F�K>��q��7��?�ϴ�'��W&7�|2de�i��Q�������4�zl��f=�]�V����|�DK���=P�]�Ȧ�;>F� ��T
1�Jr0�{%6����ˀ+��Y���8о�r�����"�����NK2+og`��UTø?[�vwp��yLw:%�#S�M��Z�}�b��u��7=�sb"CqcP�ޘ*q즙��F ���U��6���pAb7 ζ����G(۪(4�-���!�>��V�3�7�Z����z��o��6(G��acٷ��l��vS|hoF ��j�;O��	W=O��<V9,�Kn#:6-��Ʃ\���qf��t3��VI�:�3������=G6�/R�LR'�|fIc�9��g�k�l�9$�4��4P�}#�\�@�Z��ھ�4��mF��(,4�!�3+���mic	ֺ{���x�][�^���Q�f=X�Uz5�ɃzB*�~�Aa��r�_�E5L����	B� ��[ݾ,qI�z�dYz�q�,�n{���>od�-��|T��#��T(DRcr���I��8��7��Qv��B�d��i�@�([P�/��R���P�e�3=��9���k{���<��k8R剟l�"<�,�Gǈ�(˻3C�ph�2��AD�����V�8�9���{�}O��u�
G-��E�`��#:�E>|�3�~���w
�yQ��X#�r���Ma��y�9��[KA�R�	��c��2.��B�A�l�렊�ޕ��[�Wݏ�bA��H�ߦ��N�.� �y�hb�u8V�?�; 8��e����b�����HKY�DD���=����,��w�Tj�P9/����E.Ź�v7��}�a��ر�^�{:�֜�|��t%�n����vH��q��ܕ�~��n� t�D��� �O��,B���lw1 d̪�� u��=R���'M�#�m%��Pl��E6,\��������i�r�� �32��e��p���>E�rJl��ˀ�f�LLJ
@�+q�K�3A��O�7���-<�Y�cp����%�TEY��`�:����)g�A�k�[���"̯���Yw�f�"T�sH*�D{�-���H�����?����b�	
�n�P5҂�ͧ��4���Np�^x{×W�Z�L]�6X^tT[h>�Z���1P�Y�-��rt��R0��Ġ�{��ԠN	ێ�Sa�p�-kP��d��"ɕuEe$ehp�6�/r���QYʀ��:L������\��_�˕�.�aiK~Z�n����y�n)Z�t|^]�d�c�)Zmm.2�a5L����?E�P��V����sy�:�2�2�`u�^��´�#ZM䰄�)F�g֞~1���K;��j	��ٱ�����`����|�qS@���\���-+L*o*f�4.�tou�@�Uf�<���X�:,_��Uڮ;Hz0N���W�(����'AcS9�=��`9�X�[9}�v'p�C`���<�����s��G�02O�E�Y��5����.��'
�Z��"e�˯Z~2x�Cq�-����C~�a+_��L�߿���r�LX�UB�kRs��S,L������|�F�"�~��	o!/'�g鼏�v��F���|�xkE��k�|�c[{���X�D�'3� �b�z�z��cV�	���*�7?,)Dg��[K�|ǐ����� d�3,$W�;�yly(�Vy��� �}N͋�CNUy)޽�ڿ5��蜣l�+�Q�~P�X��Q,�"�-�5��/.y�5�9c+�GG����Ȃ'[+_�n(�&Ԗ�K�J�%��M3J`fh�lp�>��O	�Ud�F?��N�drуg�I����=;�L�We���{J��R������GZ�x{�Z���$�Zm���O.b�`��<4�h^0���I�l8�D���A�,�#T�����f1��o1gFЫ��D���g�c����/�nO���0�t�;�b���Q��
��T%��_8~��P���{Z�׭OIz�Wd�Ȭ�bGbV���gzKӐ��2�bc:Jri0��2�՞�\�s�e�l��ٔ�����qg����{��q�� $�o��g}�����G�wCx����}! �������+�,k{�q���ɍmkW �*,�t�����[��Y���.�{�R�k~�)���VH4�A��9��Uhb���b`*!��	`�>����ӵgm���Y�fl���J����]\�l[Vs��#�S���:6�_�"������2Ǽ{��Z�QM�;������3]d����P�R��}�KZ��-2F�;w�ĝ��IQZ�lrH_ʼ��y��Ԗ ��Ϸ��4,��UԶ��bZ�kV;�
g��b[�9�-�5��[�7Ew����"�G9y�3bY4��!z���D��~�A�@\V^-��{1}R� ����J�c�y+Lʔ�H�X��5�k{2(�(F����h�����4!A.C'lE9Q��\��e�]�l�����1Vp����م���&.!�e�GTS�&&�����L�cbW'�3j�K�d�L��ؠ���h:ʉzw��U>�Bq�L%K"UQ��1A���y.*4��!?.3|��.)Hb�N�],��"��6�����?'-�]%�p��@���,w�3�:�s �}��@��:�<T��~U�"F4��F&���$���+H3<��0g���c�{yOЯ�U��i�C;�I+?�Ls�M�k)��3�B�}��_G����Q9�h���A(G�+�\	�)�le��v��\���>@��$"���z
KX�|q=w���<	yD0��� 	;�fg�{)h&G��K�Μ �A��c��d�~ʍa��t7�
\�ڟ�oD)"�F�ѡ�A������Y�����p�:������"��Q�0�eV��v��s}m�	�t�2:���5�}�����%-�����{�=�a�&O檚zn�{1���W����D�S7��76�� �����RS�?~bT�vkjh�]b����:��w��拒� ���ض����(�Ó-+��0k�w��O�}lV%'���A��\�T�=�D��:�2&��ש�FJ4A8����FB�/!���Rch��'pjhB7�E���#�S��mNʄ��1�`C��iŀz-4頽E�_q�84:q�r�j��Gm\���㿖�� �?[0c$$�Vݤ٪�A[�j���
�0���n)��f6T��{[o���l${n�1xs���-Z>;)�9҉\��]8�{|��NI�[ ��x��B��dp5������F�)�o��������Y���4r/����}�$W���s��3�iX��J#��y�΋գ��������b���t�]��2�4\;j�
��h�'k�^J��F�$s����olT�]KCh��m���u����! ^\�gr�,���!808�_\�p�;5��&�]�u�h�%�%��l�6ˣ�-J"�F�7��*ԗ����yf�� 3�*�ڔ>�������G=�ʕ�-r�)�K;��8�;��k�AScfKN���ݲ���^e`���i�񳔯�_h�Mጢ��4�|�Z��O]!2RMbaBl8�q�j�_��6����
��|�����:|��S�l�'��lp�M�ޮ=���3�*h�6���[(J}c?C^�c�(FZ�Gr����,��r�8CJw
�B����A�5>���"��!��� w��}T�U #G��U���(�}/��8�j���N9t ����1��ⲉ��|���7�b��N,b����St�����i}�R�_�J=�<Q��y��]�����8���MHGi��D	Ī W������	|��%��wpYV�Ċ1�\3��޺e�5���>�f�����_���\n�kR�t�B�wj�9����V�9Ȝ2+)�tY}�?, JL����Dz��Q�G=��L	���^T=�Dg&\}���o�<w�J�Ҟizx�>���>�t���M�M�&��?C����6sp/)��I�����ّ������u��SN�mn�ߌݫs}6u�N��
v���o�?���=q'�1���y��m����"��W��37W�|�b��x&o���o1�M+����F%�z���p�n�d~!ct�m�O�l��Nĕ�F�Dd���g�����0�ݓ-y�|�������ttk�����<��^WX� ������X�>��r��I{nqNQN��X8x�O�xuءe"��	"�`<ĮR����"����k��0�f�h����+�0�#Ws>m(��-�}�N�7�����_�|輌o��܈M먩��+�f����f�q\��f��F��>)#�`ip�[�I��4]�-�	 ǥWG�fo�#j���J{��ƈ�����s��B>��w�&=���O�H�	E�$��S���廂L&^�<e���Ѳn�RhI�͏�;�(]�� '�t��3M�S�Ɵ��vh�A#�:i [NR��^��8R,CX	zQ�e���Դ�^l���j��}3E	%�8�G��O0	��Q��}��������@�k�JR�m�%>�a{d�<���}~�$Q�2����>� H�ɢ:��I���"
>���Ŧ�u&]J�50��Ŕ��xͲ��p�p�̆S��:'�_#>�R�����/)x��S�^����j�@�ԎS'�|R�5!S&�5�h.�@ԣ��mب�f@&�#�/��:�D!a�.7�]��bY�h�h��̙^��{������Y�3TVB�Q��>O����(�y�)�(�+�Fk�&\(z�azU��X�"�P����"�7]wl����Ԙ�����th8�K� �B;l�w�G�_$\r��0���������^�
�~�b�u�f��l�"�b�b��pyQP� z�O��/�����49������;�l>vJ˰���Cl�NH��0=���n��}�ɽ���g����d(.� �=���I������%�'�2��@�\����-|_��|g��ZY	�������b����PN��`4O?SAz>V�?��}J���!T�L��;\?͒����j���V ~��B�`V��#ރ�����!%��#R�����+!����*�j�"+�$�g�24��7��ǣ�pZ�f��'�����w�rpǳ��I��g E���ѳo'�݉@R���m�뿶�T٪nteȑw���$v(
p{���<��NB%yMj5��k2a0�R� �5<zg��N��;�&�Տ����T���M&hB�� ��y�u����n�̕N��'o�n.ÂO�<'��򚄋3>��)j���Io������p��%E����n�Y�ǥM_���N(��i$��}UbV��p���7.���g 'Ujv4�)0tM�چ�]���Z�ܼ�E��D��=,7 ��Y�A�"��O%�4M��G������-j��h��I�f{u@]M�pU/UA��L�3���4 ����d���5���j�tv$�J�{�h�r�"���F�,)��V�CQ�6#H��.�1%�E�C�9�'yl8r��s��B}P-�d�mŢU�������RrS3����٪���~c��bQz<��~-�+����뼻���4����s��|@���E������>-�ݻ��0��)̉���t�M�^��/��Xp���E��i� ���|�����T},+vT�k�R�>�Zesn(�g8e1�."<[Rm��.�ͨe��H�Ts�i�#Xu�����'.H�!����J�㬆 w�8�j�������z��7Z	'U��z�@�tE$�op����C�NI.	�f�BD�ܙPw� ��b�����,٭^ޓ������l��E3ē>C���I�U{|cNp89���3���
P	��rˁ���ŠB,R��!2�,�P*jkN���;Pg��{/�6���4@^������Y������}ҿ����H�q�b��V��#Wkɋ��� ��|�`D��"X��yP��IQnJ�}�*܄�3S<�o���v��
ܤ������usB�>�}Lnl�\7>���2ǧ�o{К`c�Ŧ� ���8���_�hu�K���]�Nt�_:���劎,qO�rp�+�����ņ��W�&�˼���4I(bB�-dh)���4����gl�Sv��~O��HT[-���ޏ4���K��y/z)vW�FI��(��
�F�t�g�G�O*4Lm8 ���+E����A�t�JnI�Z�����/�=�Q�=5U�BN���R���
h������=��==�w�w�rC	�@[�F1�A��>����L��i�k�wEiѨ��vG�����vI]���\�C�[j�?)�&P~��M����������L%Y�j�lC6��L	z���[��}⩱5���+.{I��/���Ԉ���Z�~���L��@b�I)a��O��}h��	�I����c�n��+C%H�2�n�*���O��͚�}�I66 �u�(P2���w��i���f%"�T��!�Ŵ���AiMr�C>ߛ<Q�����;��F�srF@=��GQ� �����N�/iֹ��6ב�fu�B��:�G�|�»Ԑ�X2��'���=��Ӯ��uv��.�w:����][� VJZJ��\�����hZ=�פYFN�0{��g�R0W?��Ό��QH��;1��T�m�R���?uD�]�Z���	�TV���GL��B*hf�&�g�S	^�0v����g����l-�N������˦sc�0�$0j}���E5b-.Aruq�-M�p�gn�d1`!�~N�M�;�@�}�O�Ϋq�}�>c;dcob\eG:v��_����s��� �Q :RR�(��tϸWdw��R��'����^���ş���X�ua�k_���:�m�-�<j�U�`R7w�L�BRm��q��hk�_E�cv�Y�	QV��"2�VE�5�>�t���w�Gy�*�O�� >aNq�>(;;��-d�rHS8�+�!t~RN�����&��H~.�Y��;7W��\�1������ AS�?[���A#��B�F�tkJ���2�C�V�2[_~���cF3�g�Ib�ܯx�P�jP{m��p�3<�m��Z�-RN�TVe�|�W*ĝ��rT��'�6+SU�x���S������e�q�Ѐ9;�����ۼks5�1W�㲊	����BxW���I��v{�#�qL'�?L��W��=b"��,ѻ#̃���;Y���� ��C��������Td\!3S��ƣ|�$�<�B��8xN�"z��#���ހ]��9uQP�X�g_�3���O�#��`_��K|腭��$���|łɯ��7_�_!qj � �.c�)1���7��$�� ����8dޏ_��#3:���i7�u&2=���g2�S��I�rЎ��_��>�	�=��P3;{!�j�V?מ?�c3bY����0��y��mx�"�t#��Q$��/���'k§��0�:K�]+���!|YL�d�f� �x�d���GL:�KN�[����B2O'5t����n>?Y꽸k��e�}�xdeQ C�\l�*.:��c��}����*����L'͠sTBa�����ݑ׮�S�k�^� >&#��� -��ޒ��yq�?�g��#s�6��K�I�@.TX�
q�&���.�����t�^�{ZR���<�H�i}��ft���\P�S�'�2��Eb  Q�Z�'s�5 ��i5�����G�ZR2��I�#�"8���^��h��T�\���� �P�� B��C��-T�k��F��_�}XY)���s�IT�﷛����m�?��t &�ε$�2ۓЃ\���Yze��o/0�El9Ƹ�m�Ǥ�aI��IuVja-��RE�O&`���	��
�o�$��N}�TR>�tp���ݻ��&�PL����N��W_q�8�9<G��O�����[�J$�u &0md�ERY��,����F��*����{�ZX��a'i��T�A���>��杚z�߉�����*dS�!�R��1�-,~^X�K<�W``LΧX�B�ls
�t��7�\��.j� �
C�7�\�&���N�un|�|����W:���[�F��3<v�`��%�����:����ͺ����~��b ޴�Ϣ��S�n(Im�_'7���}ꆡ6��_p2J A����h������p"X�s�c�A�r��^!� ,
�� ��,�t����ɵIO�?w'c:����X�^�e��kp2�P�a����gH�C|�U�>�1�*�	*�P5[�l�g��I_&�wb��H\�g�ؘ�������iy\�N�#��8�;&��y\��4ܶM����`.vb��SU�.�@�ړaBkrX���K�)���Ж~��(/7�owq�`w�<��N�h�<�/6<���L�"ԒeL�R_ݻ'�<6�Ѿ|*�l=�8�W�<Lv�g&cc���]���Tcr�>�lS�?qP�Ȗ<"q�ar�Jjhwvv!������@��]��(�rA,#2�O������m~9��θf�He�CC�v��� }}
�����z��\ҍL1�N �U��Ĕ�2��l��Ul/�;����Y�t mCh� 9�q�{T��J�OcW��Ԑ].&u�=HW]ϓB���9�6�\g�S棫`�	�_�j�})"yx`�L�������3���wD�1Z��I�
k�@b�Pϔ�z��vdm?#��4�5%O���-�f�vY���u�)h���#<�5K��s�����P�.3��8���C�w�NhQ���W��)�ʽ�3H嗨~��[U�D{\�o�	�3ys�	�>����f�%��؏l�q3��Pyt��d�U��P{T?���m%HL�ߵH���#0$�Lv䜹�3Aϵդ�Vh�)�ͩ�|Y3�]�����،Y��6�U�S��'UT5wӀ��ó槼A�?�GT%g:�Ϣ%6��Љ��^�F}�]�	��w�q��	i�����h�T^��\&������<��?�]ۦ]55D'�a��,�|[�\��i���)�S��L	�2��_����p���4�B�n^|�	�M	bf[�r �# �*���P�ˁ�^��&�%���p��!eQo�{z1�Y�|��}O�UG�|��<Ԃ��Œx�jJ�	*M�"���.�a�K��S�X/��ی�sD��>�Jʎ)�l�zd�kt���y6�R���|��"�?P�����dKţF �����D����������N,��ϊ��u�p@-�(I-h{M�b�2n�X[�Y/��em��u"N��W�ͰkI+�^v�S�~�k������c�Xt��VZ���y��S���6�0
sƓ��תn����Ug�b�����9Q�jOp� |2px�(����/;��K-�xZ��L��X�� ܜ�F�5�&���o�
�_��Vߩ��\2݅L�/G���&;Kچ���5W#r[)����G��igl�(h����}9i��nN<�w�8�_itf�S<�8��61��
=%��A�x�09�/y'wg)*_���E|	�ø�h��[H�~����/�|+ ��ı��@��t�("��j-�AF�Su��T���>�"�).F 7�W����$oT&��"���c�⭈�$c����y^3W/Q�OXz�Uqοb�e0��Q/����+ e�G�[�e�GS�������]A�We���mV�q�᳊.�Z�}�Q����]�m�mq��0"��1�N�P����ٱ��z�Ϥ�v�x�d ��$em@��Ѿ�|W'm��^$.�h<�T���64_U������4B��b
�b��[k��Ri~�|����ٽr�����&�QCtF��>tdn��J��--�@�/�\{�&�@��l*�eF��|�M��F��FB�~%,�w���r�eF��%�'A��^�$?�d�Ll���:�Σ�tDH<o���j�����@��ܪA�4%tܻK0�2�ZKk;!FE͙y���r���X���d*�($y6�y.
k�Ӊ"B�{W�B��腭�M�,s��w�SY&�yq��~6�coAw�u� Q4�(�! ���l���\-��O7(�l��{tpf��jl-g�緇;O�&�B@ ����@�	T5��
��r�ܩ*�],v����w�9!\�)��Ƞ82��!�d_!���^�jЙ�d:x��?]���q"D�DSw�:J����X>ZC��~=��}Iz���c/V�H�$���&��$�>�xw-4��"�L��)�4LTz~PX�tH��)r;B�>�N�T|�}"����㼽t�y�>�5�q)�H��q4��w�N.�FA�:`���� /
Y�Y����h��x��� �m����}��p_A)��(��=��"��SF:O)>��Q���0g������A쭇��;�BB*/�ޠ'�ԓw^M���}&^� �|0!�i������ [J(�a�Sx����®%�����&]?3B��E����P&jM��>!����/��8�1�.pSYjo���ꇙ�.��u���z����̄L�]�g�IΟ�����(��
���3�2M��|��m's��o����1�M�w�W��Rr��6�秖�]�ƅ
4��t��"�r��2E����C��9�z�u.V8'"�е_�� �ە,��b��К�آ� !�g�
{��6����Ő�q/#���}�@ٖn�Sn�yF�~�b�8��p�{��5Ƥ��jJ��a��xu��-Pd��%"�!! �d�O�̪�+�����`/��=��Fd��nJ����e��]of=I�g�2P��\;��o�w���������9/�S\>5�ux���foqJ��Z2�� �4�w������x%�����聭=![�������4z���h1B�ї�%��j��/�p����(̚������C�)����A��)�����l���O���z�<�Y@�w����J�9��{:�%n�2���0��_Y����eLL��N���:��"ݤ�PFN�B׽,e��a��@4�m0����ca��%;Y̹��k�'���P;ؤ[VH�(R�ޠ��D��"��礁�H�~
�1�f�k
m���oƧL�B�K��p�(-�=v�Q9����U8p˨1PƸ,m��u��R��L-tP�깬���p"� �%%��h���3�8T~��rXn�j����wB�m�N[���.�[��O4�:�]�T�� (��H�T�~��ؗsf�^���Le�6hLV���^Pՠi"�����X[�Sg�f�]@��ip�Y��3��Ճ�;�y�|�v�����Au��;�h� �E��"m5���?�����i�2�#Oj�'g��#���o�tbD3�n�!�H%�����l׬�1���w�h*�V:-��"� ��8e��^�x�`��>_��#i��/2�����̋�{$'jtrR��f;Y"<�e-��GWdvNj@�X�8�jF���L&���UA)�Į�\�F�������f�Vb�ɀ���B<��OIxA���rk?m�9�o�&2	y�)]��gu6#����M�_�H!�\Vj؀�?#����x+�p�$"0��(��B�04 1E��z�Jչ�9j��E�Q7��F��WԑR��S���M���T���|�o�Nla�f�=��Uwnzl��c�wD��`��>�M�>5���48p�r��}d�RF��z�|�ص�l�M0ۘ����
0��� "��;�ǳ�&Jȑ%����a���̴}�����A��)��}��ao�6㽥"�m��1G��s����L�����^�v���P��)��A�Q}����U���D,?^��#e��=�7���E��"J�!���xx�ZV� �������O�a�؁DCMY��<���_4�7�o�,R}�¡>Ŵ,�"~�X�0_�g�ٜ�I"��d�7�z@�ʍ�K u>��D~�ۢR }�����/V���((�An��A�h���?�u�}x�$�t��hq7��]�xb;��\��A=����[�f�X��	��n��0լ�l�z��k[
��
���8����oȗ�_�`�Fbߪ_x[��,�>�R'��S-{O�t�b�`&�1�F�/.!��Aw�:��С;7nTui���ȱ�>�����Z��h�;��f9�8�n�D1~�e�OOѩ���9��~Ӓ�S�t�����7���ON"� ��&�{S	�o�I�69NK�pkK���PZölJ�x��i&�&KX5��u�K���G�h�emgC��쾫6g,P|�喐�q��蔲���Hy��:��^֒V�Y�^ܟC��� Pe��2��7�6> URYX�M�4�.�m�د�0<߹�@1�8Ew(b��Q1NtD�2�
K0���_��/!+�j��|?o�4���R���d?L9:	�s��;HE�4YG����+u��C9���P/��p�&��� Em�	M��*��4O�4K!�^��0� ��@�(��'�(����j�r6k3�<�cJ�*�z�)$�w�	�"�ZF��yCܢ�+������L�D�+��rV�>�^�댟�l���J��\�"�e$�t�v�����f��(����2 B���5ƌR��y)�Y�"�N�x�59;E�L��@�Ͷ��aQ���
T���J#�C��G��r�i�iY�.ل�
*���a}1������"��n:m�Qb���;�q^r%�3��<�@5�-;= #��x��	:��e��A%���h�^K���a�� hW$�������7�x�{�,�����q3����D����+.M�I[�Vp��O�����p$*�آ�ǫ*)�z���>\廩E�e����M�9^e�7+_�Fm�F�a�r�ũ���b��7�2�����	�o��$�U2�� ��H�Dѯ����j��QhY�D}��IT�-�}�Z�o��2�����KDZ��^�c�$��juYJD�mvlvPl�30s[�n	L<W��3�$��%�]B�����PT�Y��C���f��E�o�IB�i@vy�~rB�b<��Y�1�"�T��������q1T�x��5�j�A�������Y�����+�p�#j&g��Nd�SOk�'���T+(x�� gL��5	��#l\�l����EYxO��:^�с����B?`�N���H�_#F/��C�S���!9��,�_j�a�-��M�I�d��jh�N�i��Ľ�����2+��~\��[��`sY���X*VX���ݶ��$P!���c"T��|�R�vKv�U��0��rҪ�-c��I'�~	#�i��N�Z7Pco@�[���k{b{��a�8�������B,�Y;ݘzF�k!����g]d�x��<jև�1$��T��g�_��G�C�k�{NoA;������p"�ڮ�J3�t
Z̿.d`t�����_��<p�@�����b�&g�(;�[��Ybm���g�b�3t�Jb%�g��L��&�;������u���X�X����F���]��<u��H�Wr8h��	��@�V|�E1�;/	����= 8r˙&��[����?>����@��$�N^�!(!�>��4}h�b$���G�SD�R��΁�ON;�d�7X7��r���焰tTh$5 ؗ��dѻ�x�����f��{�l|��o��Ҍ:��k ��� ʹ	c ��pf�hCΌ�B�k�i�]uX��k'0EJ�D�n'U	;0��"5o����>�n6e�P���fh!x�AĀ'͗r�����Ju%��@���mC��Qv������9�{��';�/ޘ��9���H�yŝ*�&+�����]�A��&���{*{��"��|�vu�o4�\X߹��w���2hU6no�۰8��4Q�c|���_1��S1"���B�V�U��L�&W�c,x^�����u�
!��,:�x�q��:7b<�z��E���S۪ׄ���\y�VE	+(�#'� m J�̜�vm;�-e���o6�̽�x�}�2��8���Z
���f���:�!��j�q5�kS��VX$s��>�
���E'v��CH4i������J�b�u�G[q����a&BX�:��j�K�6U�IxpB.��S���S�� L�g_�鷜C�!H�#Y���e�q�z"]փw��S9H`�C��K�n�>���s��;�B�E��������w3����0��H^����lg�l���z���N~X7��z��V���UQ�<��̀�s��g�BI�z�I˴zl��z{�w/�x�?�E�^l������9��5YR>T��W���K�ȫ�D�h�]����pu�Iy��d��Ŵ��˅ �k��"o�}b��%�ΐ�J�	�6)+�x�����4������D:+F����kG��A9u��q��ߑNU����a���abT�j�3\��!6tXP��3�)���鹑��tU���u:"6��mr���Uorr��ٍ���Ś_N�{�\oӿ�����k�DKk3Z����c?b�,wk�0aY�1�<��Y9�r�V�pn7
�����l�T���{G�a�o�\z�~�@����U�y�l�.x�寍`�:^K����ѹ��!W��^#Sl��1�i,�K�'Q��A���$e��M��A@&�z�xu�ͷg�aK��a��'�A��R���pڡUZ���u)h��s�+%��ܒq��mM(G�xS8�!�W9>G��<��l"���W#�O��<Õ���gU��V��>�fZ� 7��l�tgD��Y����w���̃�ծ�	�07;TA$A����u����s֊PNJ�L\�����:~!J>1.��U�ћ:��~�� �:Z�e�g��+�����zܰDS~�y=1�88��k:
@��� �W~W����|n�.�*���c|<����Jab:$�h}!ޫPBcE����T\�����R՞�p)ڥ�\nt�_�F]��+&��=��ڔlvL[�ߟ�մ;t���ye�'D��'����?��j1��?�x7ˮ���lڰ��~ V�����	�	�hp�d�]}������vU�Ա.�O2��~o����8\�M�r(��~ՓV($����� 0�M��J��N�XS�&6,�㲱�do\)�i d��߁��ì���:5�&y�yH��R���r�YI�1^T��;���M?<��eg��N�1�>�0Qs��M�ܽ����9�;_tĚ��!	�&��4�ca���;��Y˒`�gM :���O���}a�q�) X�P�A��j�I��&<�:�
�ͳ~|hS���1�X�Y,��֥O[|����m����5���2I`���]�� ����7+��\���5���}�A��X�8���Z�_�*Ŷ�QP�6i��a�%[*k��8ޅ�?�djQ�r��J'��y����6�N���{�qi�r�,��*E+��1��
F]�:�GG(�4?�kj�9.x`�V�I:�%8��El�d53rJ:݆�������Û�o���8y���)�<L	*@|eڛ�� �c�����P�i�A!�X��=��Co5���@�<�{��&@�xb�jַqo��"]�d��U�J3��mM������hQ��d�����T�ew���N��l=9y�[�a����V�E�J��#Kء�*!#.H۷�79�8�z�-���������Q�	.~<\�|�]S��ȋ�oa�ä�QJE� ���h �n��Y��Se�6�$a�1挡}F��椼m�v�lrG#(0lG�3qf�{��O�[����|Ait����|y�(d���L�Lh��]v�L%)��9$8�d���]��̝�Ǭ�>����'e&d��X��L�|s�3�(��|)&�2V4ܸ345CvN�?1�z�4qʹ�J�;b�k����Q�0�-��oְWX��N��7;Ow������!�;��O�̘�K�f���H�Y�_0�V��+�.�f��X�J�5y7�l�S����Y��HJ�R�^!�F���Q��D*Gg�4V�O�I���Pt;��N��d�Zz��(9�_�&eʉnpZBtI�2blY�Ԍf��c�UC��騂�NCe����?�Z��E�<`/�{鄑ᬌ�t�i��3l�r��ҠyV�h���ŵ�ͯ�(�IA��j�O����u�hX$�~zJ�0��v>�#`~D3�y�����#��4�n�7T��i��4�\n�$;/j:�0� 2�}[��?�}�N�Xw��avT��	� �X��������,'k���<ެ�<���g�HF|�˻�����ȋ�W��_':UO��3#�5��#Y���Z�����y��j-m��AX$o������߱�Fd�4��k�gD�c�b�Hk�#�t�`N�S[ ��!<����h�j5�]X���坐|�E�'U|�.n���hX�N�=�<�y�tT
l���e���ޞ��s���%�����&�ϛ#K��؈"[��|rC��P���eg��ep�/�8��UQ~D���k}^���<����S{�΋_��w��zo�!`ƴ�5Pz����s�(al0���\W�\UR�k�z(50C«���"���d^�zw�+���V�j4)Jz)��a�|�
�
 �����~߫9Kq\sn�e��q� <���ȧ�X���s�C]�� �׋�zR���t�)"ux�����K����ܒl~�����t�I'�?��d� Ĕ� @��03�_`�G����T��  �� �R�zL7Ǽ���^�ZW"�;eN�R�O8"64��'�lr�Ǚ^1�:�u�"����+?�:�T�)1B�L�b>W: ̠��� Rk�R���\��-��gL��9uo2/��:���,�R5x^5b��k��������X2�4�%��3�eI��CY�G�����G�֮��.>Dmf���>����)V����P��Hi�ɡ.s�LJ�A�B
�~f[9jG�d���8A�� M���}���cRx*f��σF���/ף��d�����kMɇ�H��У�[D��^jÃ/�{k��23?�`����Ld�����/�\j��iU�{��A>�c{�^�@���x��x������Jɋ�Po=�m�s��2����ۿ�T3H�G���\��|�!��$e<�lVT��� =3�`F���X�a@���n�f^D�78Ĳ��H�c��
��� $�i�ZU�d!D�Zy��+I����w�-�K�<o�~�Y�|답��9�fH��d2$�@wF��Y3�y���+����eu� M���H1�G�Z�yJ�?Ve4������~�g��T��1~���=�F��V*G���s�2�#�C�GG���1�L_�?�)�|�#SD��0>h}=6{�ޚ�RM䎛���f{Q <]�O�+ӫ؉��/Zr�'|��x2������QɋV��j�@P5ɯ�D�m����`�婚LT�<U8K��|~JDK� e hӷp4BW�{
��̜��T����]���$b�����_@��f�u��|x<M)��P��I�'����5�L��>^BNO^�9i3��u�u���
xwc~����w�&���L�O[�4�ZXy*]M|�4��h�hãO~|�;�FO���4IP���/�Cl�q�l/��������;��:-ml��dh+���!T�ㇽh�.�	Y,�f � ߜET��7��0{�����U?cڊ`�4���'׌H©�"��\�b{���Q���t|qQ�$<�;�8
S��`D?8����T3cûX�e���ο�Q������������k�J H�Î1�Bw�~� �Ͳ���L�n��1e�/R�:�S�x[9o�(vJ��1��N{��z�Z��~-b�������~�)�Pw�ӓ�J�ޔ3?ձ��Pm!ɬ��ؼ��f��t4��|���j���X�nU���&ݣ�Q�R��^6���Z���97��}ʭ�Սj�%7
T%���/��{�4&O2L��s�o?�ok��R+/��гV⇘�ew��~����,�Y�����[�0w5���-h8� ����uB�DU�ܫ�����N��������6��bV����Q�c�N-�9Y��r�����TdݐK�;�k%,���0*����9�� LS�����wX�iɫ�g�{rK9�X�!+��~�YꜺ�_xG�E�F|0\K��f-��R[2bL��8�J�l���a"gâ5[_��1og&&1��i{�� �����;.� G_o���r�=ܘ�=��h���^<u��;��~z��t��(~�	��ZG:�q�苖'�n8�>�C&#�W�~��XqK��5��
�W���1��qa�5#�왊Uh�QDXPYF�"�8sT��d��ʾ�L�}g6�B�ɞ�U�z�H�i8	���k�����#e*��|�!qQ�8�&���0�yX�}�P�(^'�w�����|F@ꝵ�*���2�ݣXo���̊gӭ\�<�/��������d4%ش�5�VX���F�8���}���ە������G-U�pQ_�G,gD��j�E}��?���<�.-ռ�dz��FGy�}�>�j/��܏>��;a��5��y���|`�R��}zUj�	ZJ`�q���;�lO�SVC��+J���f��ùjU%G ���p�L��(�������}�Z��h�T�B�G�Pe��$���A2'T�?rS0b��r�8��k���@��o��d�����}�C��������b	�ڣ�9���G0%p&顔�#`�a e4��~9a=a���bT���y� �ip��{���][����v�5�(�h߬�A�}q�)�N�-��_1O]ql(����%��9�i��Ӛf=�-���2�39Xcϋ���Xz�c
�ӥw�<3�a�����gw�Y]��sSMӷ%���3A��|*y���we7�o�!�eDL���[����x��/�d`T)��������}��b��IH$�Ju{@�!��$��%� ��fV��1�� ��<�|�1=��ǲR������PF����S����K�i��a��
������ň��AF��nK}|n���f$+;?���i���C� ��S��hAdR�4B���K�I1f�dK����"��������U�����4��9O��m�h���G�a ߂���=�.2�&(�q��赫a��<dp��|��ԙ�U�P0�Z����������o�$y�D��Su���]�b;�:XY�*����]�6)T<�j�8���]l�Q���"��Ű�����(VQS������y��T��w�',B��#�m�Q�����K��\#Y���Q���3縉�W��[�cU"]��/� ��G�)�� v�T[?m_Gʋn�Oot�՚�c�=�/6+re긹a>��$���Y91�����ķԟ��	�M����۱�Fj�c�@�GXP��(�o�D�hqf�:��aIV ����%"v�<��N�'UWV3Y)}B�s�Y��~��>��Q��,�-y!��O�$Y1ZG�F��v�	tX$��o�"�"��Z'"u@���18O�=R����F^�׍t;��f�č��kf�d:�wT�]�%e��&-..��{F�\f�Cf���U�}8���#6�ڙ?^�Z7�	)賘w�����3.�At��O| �P���SF�$�l@�Le�2	�=:�^)G�ʙ���r�Z5��A,t]��0>��_I~�R������������eI�>3÷W�3Ip�rQeS���î�4^��Ϳ9���jre�9FQ��	_lk�5�s:k�{FK�����_,B��@��%����I���_>Q�tR�~4[ϐ�� [��P?���5C:�ĵ{�Aow��:��&�N��*l=M-�s�Ώ7C�F(;E��p��ͦ|VR�瑒�CQb��E�o+�8�n~.�|f���gvE�mg�듥��KU�3<�X6���ڰ��ȿjɮ������2�]��C����W�߃�HR��0�H
�t���_�a2Q�$��E�>�3}qu�2�0[ِq���}V�����%wc5���P�`6#ի�/*��v�`��;��ǬL�S�?�Քj*R]�aȖ�] �� ��j=/�����*��C&�D~���PiK#�ޙy����<rx�y�:U���*�-�̵$�!,�*!X ���a�.w�G@�]��nS|�B��H/eߛi�X,�uh�v䟔$��߸.g�l�G�k끽.���	�����ë�?3oд�؉Jz���f�w0��W~�wz��s
 ���6gY~=���L��f��Jԑ�{ ��y�L�3$8E�"��|v,���tW�W���Գ8^����-�T��Hx]�yk�J[| �c?���R}�=���~)�8���gUwX�c1<B)*_�cɽɱ��{��
�EGf���I�L��V���k��bn���*��_5�g?)@�	�c)も@} ng'M#j����]���݀I�
8�C����QYߖ�3��W�r�!ʮ�3���E�E��0`�t�ju�pW�^WM��[��xI'T?gK�j���G��:jm0.v0�z�\~�Ax��y��2%j�q�Cq�5�A���F�uk�}gx&����R^*����A���C�I���D�,���2����ϊ;�0�w]�}�w.�^4�N��3��-�n��X�c����#E���!>�d򅃲Gu�&n��K�٨
<o����L虦Y������D�)�3qM"+�0�)�w���[;�'�T0b�\��F��T3�2^��A���=3FQ�F��JC�[ᰱ{�B����n՛�c��/��9
�'>% ��2�!���P_��5�G��[�9�O�i]"�q��_M���`��#~Ӝ�F}2kf����S�92���xT��B�
�p��C�����W�򽰑�����=i�ΐU�$�^�e(��u����T��J���M㯌�o�x�ؗGy7-Tѵ2ݛ$^���Yy����_�x[fq��������N+��pN\a�j�S&��c;�8|S���?�������`��x���hA�����V��ۨ��;Ic��$ ocK����l��7�I�
�M��έB�g馭O�]�K̰��;6��S�B�����g�N��YC����[�m^+4l��@�9������ �.�VYF�2>ۂ����tg����Y�l/S���+zHٽڱŎ�"�y��ڧ1�^QT�a~�Cud�R�XE���]����Y�H�|*	+�(i�Jt+�Y;�t�8Vsl��
���q��6ۺG�B��F���:L��Ad��}���n��^,���m�`��������:B3q�P�}Ԩ�`����x��BT!�+�0��t�oxH�1�i$���9������/�y$��'*�hwӸ��\��L��ҳ��
s�Fo�m����WZA��S���<�SZ+Z6����nf)�������2,��'�ӾAd � �2O ���Cc}�T_إ@z���k�B��H�����AA�t��lM|��*�ϟ�d8#�|�D�b}>+j)%(�.K���4��ËA����`)��F�dXX�Fy�R�X��l�.�J@�R���0�
�F��}��*���S�ٜ*Kz��`�,�t^�@�)(Fq����F՘�2��!:+���}4�F���ѯt�]���[zi�����u�T�g�Nc�c'�4!����9�dJ�b��FV�)����K�wd~��5@��s�"J�1oI�	|F>ZDt�����IX�Tk�d����O�T�ڻ�X3!� !��`����ۇ���p�n�&�F�f	�L:�f?+fJG�����R7�C��
�c�g�������'dB ��Q}�ww�k/0�р�TU��6x��U���rw)�Ba����dt�6���^��N�"A�}�E�d�CX���'.:��&�7��\:��&���U3����2��1?/9�Z
����n���ͭ�ڛ������eq�������[�-����$�ri��k{:D͒�f��I��X��f��_3���oF>:9�j~'I/�iK4@���.v"l��o��.g��(�B�_Ǻ{�а$����k����!5��<����wb��*��9Q�SR����!U�����$�����4O��w�t��@�4hp�wp�:uaڮ�����Z�m�t��*7?C%��#�s�9�#>�o� �f<��ɬ�B�A�ާw|�vU!��7��y\4Nn��&�m9n�µ����o� ����9?���_3�T�pH���& �!B �T�ek��t���-!�QET��]b�8��ً�pCe�>Lə��)�I0r4 ��edv���^߻���<�Y�`::�E^�K�
�G �ǐ����ý�]MպyNm�f��p���*R 2�8q�T,?m�vҜ-���2(�3=���57k+I8��#�;.���6{D�حT��U�����y�E���O%-� �&�C��@>����c��J&��m�|��}k?��N�0�$L+`���w��s����}[� �rՆ�PX��l8�3lx@z�l�t6ad�-���d�O X�\��1�M͹ػIBM�q��0"�ޢ1�v.nҽl:̿��"�a��u����o��2��� �u!*�s��^Ԡ����~�k
�w����⚫#<(/Ą_�Է���k�kJ��]]!{%Z�f<�G��� u�+�ZbrM�������gtI�ģ4���,W��e*��|]c2�I:�\��5��
�Pѩq�o�|�u��5��81L"Z򫰈����/["#��9=a3� �1 ^�F�ͺ��lPr`�nn�z��_K?�ֲ���WĖ���o�2���_^F����gVu��@�	�F�CX����GJ��ƒV����r�o���]|S&��гt�n /Ś�|c� mp#��'~�4��R4i<0����<23k�������֝d��bH4��6DY�7W�S�|Yxo�ڶ�g��
���xb�nW�qȋ�V!p�Y1�E�2yV1@�/j`��Q�F���A�B��@�#v�_F�H�٨6x�@�R��-v^ܢ>�����H�J��@�}Dµ��K�z>����p�jT$~��o��|H�3�A��-�(��1�xZ��!C�yP{^�P�>�
�F���#MT	�M1�@LD��nqeV���{ :eU���k���}��H�"�?Ik��[b:��S��z�=1V(�D=���/��'iT�f̞*��V���1,β���ۢs�r׮վr��X�_Ī�RH]�#ڃe�L=�ʚ��j<��Mٗ���[uV,�M#f�+ѕ�)E_������w�v�Pl��[dF�(�����O	7���]�L8�`��Ám�A�����/�Sl���Qa+'�IZǄza�_����&uw$]�1qW8{�l/j�epϡC���a�]�&^�5M��VV��p�`�(1�sI�5���⭚�hFɇ|��xd��gc�:�Q۫9i���P�Q<u`Q�IeQw3e	/0k���X��CI­�A:3אּ��R����ob>̬���`�@����!�Jq��g
W-<H�ڙM��V+��bA�D;�K��`2W>��=.���W�a��_*E=���u��lu�x�'H�u�{�5�:������pq��.,S�G��"*�v�ۨىh�]"ͤq�(�z�>"w�I���dN[�]�a)�U��o����f?$��q�BeM]�SW�e�Wy���RL��g*�]�*����p�v��c �-���qK�@�����F��*�5�J
�&�8UX)��N�(w`���+�\2![s���[�ٙ�XJK��%n Q��ң�ϣ	.�W��=�����^�RP�A����do����"ڭ�g�(>U��yp�ר,��A�0��g���\�7-S֤:g�f5�_�5sf��~�[o�0C�@�)�3�/���*�u��TD:T8��N��K�1�2�����ʢ���X��6�z����X�C2�b�n�,��s""�-��Y�Ԟ�+CQ /�Ux���n=��:��ڡ�F�-�y#q~��b�{xI��k�k!,�,�!c�I�����u�,.��b��������	�Ҝ�����}j�$��yF�ވyX���\�c�V�d`ym#:�5,R�����7P7p�]C�]�H���0<�9��a�xDf@g����-���l�@eHa	8|���<F>��mz:�}�8��/`hC�`G�1u[�@1�� �1�Uz#��:�y������A��q,ҲR�d�q��B�͉�>g�n�P%�y6������{%O�������J8�J�7:�X�A ��b�}�J�f����k�x!���,I����_	t?S0
�^pݖ��$"����L�q �M0��Ϣ�E�����p6>L���H�>hH� ��ђ�	�Exo�KY!gm(@M�
k�'~I��g.�JtɗK,g?���apv>� �pР�����q�Y������e*h�	�C���'BM	�����7��Vo]����b!����)9/T�o��qSC��P���YLf��Sj��{�	M����+��H��F7�d�!V�3����Np��B\���;N���K7O3LCj������M۽I���<I� {�r�ޯ8�3��s�g5+���i�i4�x��!ى� ��u]��;ns#]❄4��S��;-�K�j���v������n;;�<�ݟ�V��������v�=�G	�"��<�jz4s
#�E�����\?�蟯�ԥܱð�� F���6��WM�n9�~�u8��i�ܙ��3eW��]*�Ns�jge�U��8�%�������-�u�ȶ{i;:�O�`'��&WBv�M�F�q�ߊ[�.�vI������Z����ME����.yߡ�N��
�y�Q>��<��.���"�����7�GZe[��&�`8#R$����2����燴�H̲Л� �ː{�.�pEa� ��+�9i��c�xR6J�ony+��c�O"`le�@��F�|�t3퍹@��!}'"���W������u�tP)��^$w/4�z%<XU���=�(�J��\�G�Nh[I��d��e
�"�A�l<��}&y�����6Xs��_-޼�L8cK����*�T���0��������|>��o#��m���a@�v|�4�K���b�Ko�[��w�K�f��RH��v��e���e�%}��'� �p���:�1���Ic;l!����w�s��2 �._�<n}�����M8��)tg���w���3���
ex�G�2���G�:V��4�S�y�آ����~�\Iv�5d�ݧ���M�۬�[P��f���u�d�5�*� �0��y;��_�lG����o�?���n�V+�8�z���\�^ã�ƣظ��g�%8�NY6ḍu��AH�V,d�)�����-���P��:t������L��x�2 ��∈�=y��bP�^���	� CF��9W�i[����K��Ԡ��O.�Qx։�tT��������s�l ?�S� ���t��V94)�/H�yf��@�Bn��e�L�FOB���oɈ��3H!D��a�"��%$��I��f-	:f��I�ś��֟l3BY?��c/��ϸeӫMB�c�i��)��J����k@��L�<���׌D���km�^v�B>��5��'�� �l
H���yY�y f�&�����W.,���N|��@F������uS_VG&![�X���"!���y��Cm?%N+Ii��k`RY�@���A0.Y_$����K�5����[��]=)P$+bL�Gs3���v�F�<dU3��"{#$9o����0�Ե?>Ip��? ��:���z�\�\~̗�Ō��K�`pt>�|*��"7�p�s�&9=�9��wnw_Y+�����0
�y�$E���^�M|���+T�H�7�um� ��\�����&\T��GxVa����N�̄�θ9��;���]%H}Q��{�����X@�^f�OTXL�!7���[XS��Q��.����l��U���/F�`$]u#<�e_�g�z�.�)��W�j���߉��4��~5�&,�$҇�m�O��I^��Z�1��WRCx�1F�\�#P�c�u%�K��.Ҋb���J���ѠiïB��@G��Q�ٜ�P,�=z>�6"G�g^�/*I&j�*l��E�c����`0�x��\�4�*>��
}���p����;��5v��6���y�B�z��>���~)�iI�NCB�
Wmp��ڬ��AO�ّ��E�8D�0n<���T]V����aɜ�][~A�]���tO�0P��r��:5�%����r�Ҭ�4�����ZBH�n��s�G �Ǹ�����>:Y����p�9\���D ����G�e��$��f��cI�B�y�39�Х��V�BT�9������Wc?��v^���Q?ŵ<{�b�ď�dK��$W,��CMPrVП���',�{�:\.��0މx�)�$+[ Mk�N8��`����!�@N���2T[��cU6S�`�c�y�� eF�5���tj4��H.��C]��#�y	
���\��m@�`3��	��_Zܳ��	>�ٻ���������)k� '4���0�u�f��W�C��}q5YJ[�5A50��ء[C��Ѹ�W�jy{;�/�|+�h��h9���O.�@c���Zt'\�v��0�{���2c�X���>�;΋f�>��|-~�������836P@+�6jUr�(<Ŋ�sy��.t�|�O)��~�3�u�Kb�u���֍H�����O�n�(T�^��,�	X�ث�/)T+Z�TGD����� L���>��[`��?ڐ��Ufa�8aIN��t���Lqa4���NHS̄D(M��2Wt�I��k��G�5��yB�7�3��O9��$�,����mQ������ź��{--����0!N[����D�M��T2�!�\L3k�\��4}�lTϩ�l9�f}\��1�0���A1i�LA�^�7J�s�4	1�o����r�"��>��iժ'���mrO8Ħ�P]!��5;���_��L1[�h�81=}ؕO���}��bKbV����C�qI�ǇC;�!!�I�K5ai~Q���$�X*D֤���5�!Wy�Z�KߵJ�L|a\��H�,o�9s��,ĽĬ�p��d���H���0�1�*���퓶sF�J�:���XBc��k����E�B��t����$C}���^��Y�F�vweRk���:mf�%���g�
��N_"�La��b�<@�o�X�¢����o���}٤6-2[&��3J75{g�Ka�l���4'LW���V�Ә��wxN�sfq��C���d�\zN���̏�\ς$_D+V(0.�,�0~]5;*��ӓµ�H���<yMOy���h�=����{'E7s]u�`@P�?�ri�j{v�t��$�
��9�|$8�k`YBh1�u����2����AI6��&ǕA}1S 22�n����t׽?��H"�<ٟs�#1C��Ы���kS�S#�L߿:��H"j�~{��y�	�S��@�Y���.7�fh'7.�����|��	�r��Jɩ�4���l�d%�2O,��
�XU��*iU�ț;)��!��)J�P�ߗ��"��h˟+�u��W�}�>�P�J�!�v.�dhuqb���r;�Z\�e���ai?{�{�X�n��8�(c*��+�>doj���#PeL��b*�`+9m�$]�N[�&�S�M�dCjEۮ�����u�����ri��s/�~k1��cj����FYQ��-d^q���N<��``Rp?~=��'��[o�Ԭ�����iΉ3��A���,s��1N�N����M20�^���l�!�DfGcy>�n ��'����[�>s�\S����]��K��M����W8��o|�|���n3@�[�C��]w=\s����+��G�9q�O�����8�LL�TyjGX��e�Ղ�Z��J���kJ���}[T! ��Ś�}�5�Qg���"�R?:��!��G��|�.J&O�#���ş�r,��{�ҠA�+t�J�r��V}�9oKfۥ�4`H�Zu�������#��5M���}U�+�*2L�1ʵ���{��I� ��=j��R���*a���8�m@Y�(���}�c�"r�X|�d�f�Sb�Z%��: '�)ۘ������`����DR�Y#T�inDlzv
���+��v,~�{�&��kJh���ab��-�8+��p�q���xKiebԡ��M��̂��e��^��Ѣ�1wA$C�;�Y=����ד�/�۩`�I�()`����1)�^0�� B���#��OKϓ�3ȉ��4'q���5�"�F�&��+˶�~@U.P}�_���˷;ȚN:�& 
_(��D��B�v�V�F���u�Ba}"�����k�V�f~gQ��VoM5\�0��|!��"	����F���1�Z�D�6v��ɷ��tC5���a�!H�I��-�� �y��S��I!�X%~�	Oqw`�T�l��>RF�k.<�=��jtΖ�2�|�p�<��,aN��g�o��<�d�B"�<�b=��зV� Nٱ��ܲ����b`_؇8�2b!�}�5#���tuV��z�=�I4n���ۘȹ���������ͼ�@�6�4y�c�i�f�>z(����>��*�-"$�s��X_�"��V��N�Q���M9X�ڱ�?�i�b���<`5��u���z�!u�?.sUh����)ɸ�e��(
�����9c5��J$w��#�`'$���Tϐ��8k�vRUf�����>�u#6;�auX�9��[�rX��� ߴyB�ߒK���[�̖i�s��&>9
�c4�<���0\�#. Xm�z������F$R�a����{8'�NOV�w�Y&��^~�QK�Vq��L�#C������σ*6<yi�;��3�В��n�cc�;����|]����t�܏t�q��$i<Wv��V0}��|����S�[�-&$��4}���_,�I�%�@1�GHL��ĩ4Ѿ��{y���@��� a�D%�<��H�|8�BUl?ެ�B���W��-Ca��\�hWj�*/��ce|����jy��bٜp�G���B����)�t'�>o %uЕťn���) 6�cTɻVM�����e�PӋ}��}�d�p<�I�JG&$w�9"k�]�zE�W4=�*|�Jizš�bE����ΣL`���&J������	5g�ZPL��7C�D� ;��ev����"d"����7�=t�3p���B��a:����c�dHHP��H��4ri�M9�J��G���C�RP����JJ
��)��@�fgԉm�Y�.�	�Վ4�b�>=�آ]c���7�w��]b�ՙo��E󹈆�y4{�6�8(��!� �;�����]�;�U��"z���U�刷$9.�I��sK�}�GD�lų5�l6�#+����ɻV\,-bq[hjZ�G������Z�|pNM���"�\~h������q�T�31m��Vk7Qf�l܁��*<�t�;�1��Ee,�D�
Ad�7��J�aK�U��W��l�b�w�Tg)=o��}�;G�y���0���#�����N�'�8�3�w��%a�X�y��X��*pݻKR|�;���JԹ�݌#�6��«	�[xd�P�JT��H�)ҁ�X�J�����^�qX���=�v`�Y�s����)��濉�������n��\a��O3���d�#����k�wOX0�J�܊c˫8U��hh��Â_h�*���֢��Z�s���%����l����;�*ʭ�Z#��;>�̛ݫ�5A��r�j�=��~��� w���a<Qd��J�pL ���#'���M�aӄ��H�6�> ��8ՎȣOӚ�ґ��5��1| ��J���vhW,6���PY� NS�y���Ǯg|�?i&f$�}d�S�3�md�ғP�[�Aj\f�B�Xg>ޒ  Y�P�*4�?�>��z���VݮxX��l��t�[u�z~VIt-�o��k�X�6� ����>�B���2�����1��	1="O9đ��~�T�|��恇ä@���<3Z��h�B�χ�oAK��9|Pʾ�I��]r��O2�`a�H��/�lȴ�X�0���D/�3�ߺ���&u�C-��r's���������6��
�Z,]���6	�䃝 9�qf���8�q�zd�S(;[V�����8f���'�aMʦ�:�4�S�AHR99		��VDz�s��J�Kf�:/sC�~�gV��d�M���U�ݣ~��a#���C���u_��s������b��ਵ�cۊ�)�yqY 1���^�;��MO�������
ʩ����n>��
jEߣ}%���p�Q���]��q(4{�pIs��7��{���w��3[#�휁?/�H���]4�����G��׭�<V���(��&x %�y�r
�i�ͽ�	aw�1�j�Ñl���t�2���5�.Q�fn���޲:�E����X��vy�Y�J��@"�We���t`���3��KU�Wv(���\�ߚV"3β��UV�í�F�E"��P��'T/�#��2*6)�uv�x��SM'��}В�}��}�e�:D,�v;&KC��@K2���t�|���J�v.z��4y �zu��J�3���@���%=o)�/��f3]K����jz�l��U�9&��D�e���G|3�鸈B�����6�v�>�<Lkĭh�wx�0�{�m<�_���W�Cg?�`)��7���`��l� ���w61�tŔ��W�|.tʹ�0a�4]�(9T�lCs���O� ���"X�j�!���ڴ0�lܲ/�댷�����	�ᚊϞ�[�`9�؟�JD����y�t�N!��cҀoL�8uV� �Tߛp�����e�έ�Q��P�R5O��c�2�iK���6��/��U}��7�j�M���)� �9�@G)փ\�_v7 ��66ЙR�K��Q2��:	�Q�!�;&�T��.-��N�׬��T�#��Y�P���U�yQ���b��%p��� vzْ�!>Y��>7V��A�TT��ϤSr�
O�?qj�����@�rj5���i#��Ѹݺ�>�[��f-%_#[���6\��Ld�4?�t��rL�&vڻqPD�jv5#_���vg�Y��;�(�[n �7��lbY/��S�z=�3M�+��7wr ��rv1i��`�l�u�5����pUҝ0-7\FշA�K�̑Y�oTܴ�T���
=~�M�{�%�ު�����
��n��Gl"��@� �V�K�zTϯʪd
Y�k�N�Ƀ�ʑA5���[��I��'8�sb�r�oЌ�/�8(�IT�z�"�5W��C�@j��'Z���^�v�|��k���xU�׌"?�8�R��Wf�׾�gJk��.��勋�g����P�:��a�6����9ڣ4�+jb.��Z��K1�4��Qr0PqI����,*0s0�8���9����6�����S�P<�E�;c>���ĥl�?/л�D8�E��ξ�@�$�=�Q>���t���I��ux�5�q��� ��+� /2(�����2�Y �w��~R��w��y�D�ϰ�=�
2 ��i���|�l���P���,Y\�*�����l���`�ƍP��L�9� ��Ϊ� �·��P%;�P���^���
H`r���	�
Kx�1���k%��vk� RD{w��%s�B�y�oWE��n��3��{εw��@+�-h�ʭ��:�7�-�%q��:�Wi��'I�-���ʽ�q��<}�$���n`�ћYA�����u�ƵDX�హ����lCy���y��� ƗI�"L�tR���My�0f�j��*u�Pt��~���e8ʁv�ͱ3VX�\�l�G֒�6���`��p����,+��V!��U��գ�"��&#�,:�) ��
�r���e,��+�p��J���~zcH��ij��Ox�ܼ:��Fؙ�R�6[�|�Za���cSK�Z�Ev�%S��y?vܯ��h��#Z޶UI~ɭr��g���䟠�#�,�Yi;�y���$]L^:��sDT,�u2�����B�&����RI���4���=嵐(F�����j*�,�0NV���$��;�n¸o�do��;6FUI�ȅ�L�%L��&ٲ�箼v�����"Q��*D�SN������?�����skL�s��W�<�|����
rԀb��̇��/郧S;�Q,3�*!a�Du�Ř��D-���[rH�����5RP]���xp	O*:Yx���Q��p=��|�k��!;mN^X"��\��*Ա��o�k4�:*��ȝ�7�"�~$f���;�۵�q��w�5�"��Zt�{k-�E�^ك
 ��Ʒ���c��,�N���ep������u9��:QES�ݠ���ܲ5��A��0*�ĺ�x����q=�a�[f�����.��?�@�����m�������_�qW�~�`jI�p�+���i0X�4�Kݡ�=�of�h=/��k��:�V�Ƨ����;l����O8�
���'� X�K>���G?}�z(�����`n��A�s��3����!�e!ą�{z�eH/[�oS���
�n�G��ie�3$���G{��uR�ɽ��`�_)P�;踤ȸ����؅u�D����U�C�,���j�8.O��-�i��@!��"����]*�,��*��0WC낤nb��0* P/�b@��,��vP�<�zعZhי�ߵ��CŇ�X�D�tn��]2do��N0��
�m�/�mnKe4=�eN�-zu
�����_�����?��c����
WJ1�v߇¯���J�`��Rp���euC㰏Uٵ?ifo�b�\�\:��]�G�{���0��l�'��]�����+k��1�(�KD8Ǻ������r<8yҔ�F}�@V7�0�M��b�nz�i�-js	��3�ײ�[T�F� +��&Ŗ����*̎ユ�
�N��К��U3n�f�΢M}[�]�4{��-8v��^Fx�a��ӳ=zΧkΓ^Y��ᨥ�yh�8�s��#!N��g=5[wQ�݄*���a
a27����p$�}��̫8�ř��9I,��T�ʧ�o�vsb�ۭ�ɮm�%Czf��¨"*f�0m� 	bZ��"��^����v���Q��i�a�*�,m��Kğ��q3P����������ɍ��R��B�3�F�}�ċ�/վlߒh�WG�S�֨�1��ئv�
�ẩ9gqۭ(j��Z�D�Jz �|٧�Fmq��ǳac5!����G\�St4m��<(�Ql�c�w���_5R]?�kT����yy
�؛�wψ��n��z\�A��H����	[����fi������"f�LVHFKs�
c��"�h�NV/����&��T^�����~B����Wm0{�;zgZ�S����ͮ��[s�cJ��
6�Y��IMw�p�+M̆�`�f�5Kɇ\.#k>��jѥ��o��xjЙWxJ��� �5Q\��I5~��5%��6�޹�K9h学�oLN��t3� ��<?���bAC��݇Q	�ho�"�	
8���d�'�4<�U����@�0���>C���s��A�\*��VF��ؤCɯd�V:�΂2PJts� :�\�ά�~$kaF.��y
�7�@	�5���U1��Z"�e�E�Ҭžom/ځ����[�q�M�����cOK��&��(֏�Hޞ��0s9h]Mfn\&����|vޞ�y��>Q�0�,�-)��5v�)��G���js��9��^��h��b�;�O�w���rp�x)��AD p�1�)�,d�]]eTӎA7<��#��� �}nɖa�^��2�g}�d6��_�i�~O��޼$��U�n� [̴���M,�42���`]�^$*�n�"(Kf�����o�N���󧣧)Y|�-A�^|���!��X�b���dUd5��M��-PI�o8He�pa ˺b��-��R�H8�����ˁ�+mֳ$�^�lj�nE���o�+~�����������f4a�����Q��g?%�n+0~�^%5��h�����3]�T�S�0�(��@����4�D�1׻�:5K_u���X�CG��9|ˡ�;�x���h{���>�AxC�j,Z�|�M2�+t?���e�~Iumf-WryA�l�#wֹ�p�U�45��ڳk�w����/����7�J�7��W��X���g�N
���j�����]�e�<)�D/ �����E���/��L��ɀNg��\ˌkX�z<�*�����5��o��)cW�*ٳ�#w������鉊��v�<U��fP(�=�FC���E�ۺ0��5 h�J�x�6}sT�L�W��;��##�����:1�em�%|&1�_�s�g4�/5�d����j8T�1����� ꎙ�Z��Y[��V�)�� �S�5y�T�	���TF�>�;Dh2»[��+t/�|M���K��M�VX�xV�j�38����UE���d�
��4nm�Q�q�/�mC?�uq��U*����x�b�J`���4N�n�c�)"�(F���&��@�����j>�!@ eg�^d����!�I��U���];XZ:��I����Ѣ�b��7�dP�N�۹�4��ٛ��(	�$���z��F��|�r���$��_�����Ci�V}S-�@�K,����hy'U$�4� �rӝX|z�¤�BNF�:�^8O��ԭ�[Ţ5�tL����q��B��������W̹h�'�ki$�����.$1�o��@���ܶ��n�� �-���]���L���>qG�H܏�ʗ����n<i�e�֗�]���?���Ӭ�\~����*�rM�,���In��JJ�9Y�~����H�%:��� �gcU�߫���`Xu����R�R9)
m�W�0QXl�)�n{�������ɑ���݅�C��J ܊j� v��q�m��������!�(�H����j*/C隢"eЪs��b.��!�D������4��*�U����$�ɗ��-�[5ӏr�)#x[�x��e��q���p �O=��"�G4���b�zM������zm�%�
_ܩ_\ q��Y�1�@fᝂ�Z����}��Vپ,���:�)$$]Œ�c�8�7ኞ̥y�H�C����<�������gu�X�P����)�D��C僱�%����E]b��/��Q6E{7�a������۽�Fz�"��i�Q84��#M�8�4�	�� >�Th�����ۑ������w��}\L�@�O��y[���-oK��{��1�R��+u���5�Г����q��R��΅-��ܸ _vٷ'��)tf�
 ��wZ��;�d]q0��}T-O��y��� J@չ˝�_\6y_�[3b�l,\�k�e�T@�vD�3�o1L�YI)�6L���h�zJ���ݥu�O����$2#�G����u�:�4��#�&Xl���!�-��X��5_إ����J�P��Aȶ�i�s�x��T���z3.�_ȥ�!�����6�w)Hc�W�����J K�ٟ�4��C�ĳ�˶7�ln�
� ���]��B\2�"�ԫ�V'��	���V����
�Ū=t����~����!"��(�H�%�E�0!!jK3�0:��d�^�ޑ���G.��M�KhS6�X�mP�H�Z�g�Bss���� Ui΍#L?E�ҙ �6[���ݦ�2+֧�:�-��O2�R���5!9M�@�Am�"I)�����մ�tw]%����Vަl�Mz�f�M�ܧv�Q-�rNo#M�`V��F�}/��S`��O�TK:��g9��큙�t��ܛ��sj��ta\���|[2Rq%��ƪ�U2q?�V�W�!<�Z�*1�EZa�^�pk&��6n�7Gw"��EXr9�
��?�t�\"�ù��++����Z�	��),*eD�����9����b���t�C��e���@G�sq�Ֆly�*���^u�$�'"��W,;W|7���9@�����2��n�"wI�R�|��&�F�s�NW��ϵi�qM�%RҶ�nAdt�+gF~���w�1�g9�k�!�$�Eo��a/ſ����1?��8B�Vl�KL�xKQ�]��gݐ<;�f������ױry��ߡOJ�#Lx�XG<<����?�V���P�O_��=[:j���5����g�K}C/�4*�g~ү�P�%T"g��&G�:υX�|����Yf�>zƺk�S+ؾF��=��y���`4S�8�)OQ����e�9-�H��<�RZ*�k���5���)Λ����]qAa�����^uM�����6M��HM|G���Ms���73��>c��%�̎��|��Z1���aƄ��
U�����nR��!��ߋzF'��]�%d�a�bLS�|Q�,���zOa"�z1�9������������KM�g�M��toY�djt+R�cIPe�SHCM��@���5����Ʉs{S5�I97F�$�^7�I�(���㭝�Na2<rq�&�^3�V���I��p@©�pNL{�>�)���_�X��)޽h�¡0��ܐ��\$�qA2v@�_��SQ,�LZ�a�^⡷�ndoCu���dݖ�sh�Q`<
�=n�[0�zފv����V(�W��h;��V1�&������T�Ft���2〷D�Y2Y�0��:m���*˘���&�w�l�~x>��i*�yB�2�Abr/���f�L[� �\���I.��?b�I��=@�;���DpRX�W��s �E����ͪr�W���j���kE�8d�	Q�8S�5tq��Z?8�a;O3�]CEn9�3��ɂ�2�c��r
oF��>���"P[�r,�7��I0���WP�M�T:���9q�xN5B�}沆�LK����j�x䝜�Mh�.�F�b�]�	�x�'O��م Y?�(�X�<� �`������F�����YRY��pF��a4�uX�Zw�����=8l,�x��e��`��'L-��v��i�ɇ��v�;�2�h�emi�Cl�oD(�S8(��a�����6q��E�ĲJܴ��Tl��l�b˴��L9�����Ȼ��P�i�d��P�Ve �J���¨����2��d�P�K{��P���#(r�,�`x�̞�K�cp��qv���G��VOS���IM��jLR�/n\�� ʧ��I�K݇�GN5��9-�`G��r9�NI�|B�u�`h�n���.�Nz)l�|J96�upi��G��_��G�3�y�̥
���U�2֩���K.���ʧ�M�S�Q��'��o�	[�_��n��Tn^#���*4����P�4�gwS�J%mZpb\����Py����є7�5��?��+	��tO���.��~��n=��x��>�¦�̄��`Y5:+܄�1�;�Y�g���l�/�w�t��-���ܚp� �G޿b��Q���v^��JrW `�fC���d,f���?��� ���cI9�L�U�y�t���P%�G�@���sJ1��s�"vUgy��cQ��s�fJ�Y��^[�D�i��ڟ�+�ȓ-�����KݨG���&��׷�9���^ޡ���HU K����2:I���W;���/;@&���`&:�Oz��q�y��u��>�G�'��:�@0�E^+�E����p	֎�E5ڀ�.�ҟ�O%㗀abn�k�>�b�R@<��O��i�9��,�Һ�.|k�ǜ6��R�3�,t��u��J�eO��8i.�;�x�]��}S�H���Lp���q{kBv�Kb��7�	iPW0��)�����)�Y���ȲC�h]�?�l��?����P����Z��KV��Q�˹I(�#`f���2l�'���gd�m���"�Zo+:p���YZ9��)�I[����[�����l�IE�M�ܩ�%���ʷEeiƚ~p��hq XN���muKAߏ4+�B����<2�����oz����jdTɭ���������'2R���Wf�p�x'&-pxRDW�k�E�]��B r"nj�B."�b@�R� 81�7[3vwS��Y=�|�N���Bx�:	)�1����y�{�eX��]�܊�������eV��"Thtx�	f�:���vH�����g�X$:$T=j�sA�GG^�3�+^�~m���E���2���'Ǣ�[V֗��q#�<:��5�yD����ܮ��oR���71���
�W�3�J<UpPǩ�q�Z�i�[+q^w���v�>^ah0C��n�IG�]g�✗f9݂[��l���yi�U�3N\Ɍ�+yUvBZi3�Rk����њG�]y�.�n�����-��s���_� ��S*��a�kCó=�2-�������D�l+���45��@�lܖ�R[��� }E���S���l�Ly�7�Xh�y1�e:
$F1(GU��A@$�{����^�?3�md���*ed��+*P@_�J��G�=sOs;,��ݩ�=բ&���A�d��Pr
���I?]��N�7�2k7�^�?\
��cms#\����|�u�Z��AzE�I�V��muq���J5�Iwi;s���)�J)�
�I�����GN��u�#�o��~�l>����&����b��x|�X�b��U�I�o�n�?Aw��a�W������\�,�u߼2ǅ 3�=�"�����h*����1��րyI���q��5��I�5?#���C�'$S�gS��D��������5 ���o�g|��g��R�g\c����]����w���J���"@�]�I�Ym�� �y �<4z�6���tOy_�8c��N�g��={��/b����RaN��D�����d���(�XR�HbP�O�%�u>m��Y�<Ѷ>s���((�g7�7[X��/˺y��s�#��l�쥂����	Ӌ�7�����o����i�{I[N��m
��5m�K�W�駉^�;��d����N�F����}�`f��9�m�i����$F�KY���8:�4Ԉ{�:��&��9I��.0��UwvKQ�ܬٛo%F�#s$̊!�v����cws�+_/NW���^@U�	�B'9V��Q
툼���#�CD��C�b�a��'b���=��D�m����`����Èr���	u͒����F)ez��d9�P�<��$~�Rf&�'���sZ�>$I����[�#N+c�%֍��6�_	���c���YAJ���'��it�^!"-�v��yN����1ASE�-���r���F[��!
��#��
�'؇b��s5h}��*�[�)���w?Bc �a��y?�E���b����5�nx�^��ԀLM^�]��S�P��M���
iV�{,4���?-
����,�_K�TVZY]j��`c�=����~��#I�^>���xz��\>���<�x���{��
� }x�\��i���+ݼh]�YK]�P�g�u!����7�W�+�03֙{Ҿ�Gѐ���z��p�l��������w�J��ġ����"��)H���޸o�~�ߤl�R��.Ǟ>@��i��b���3/�h:R7��Z"kFz���ԏN�[��!�F,j��3e������VhÊ>e�>�Hh�6����=yg��qO8�mV��L�dha�>D�Q:{��bɟ�_� [�O���L����P�6�T<�����:+���iq�|����SU���*�O�ZnW��d#+��W�Y�
��n������Pѡ9��b���ު��S
\O��P ���;�xz���,ުy�s���AL�!�4��?��ؐ�s�w'�	: >�l��Fq]{k�"S��]��2^+5S������@v���]�1�  ��H-��t_��7�l�tI2uQ�.DO�k��H˛�pʯz���ĥ��h/ϕ�C�o��g�4���C`&�Ω��a��{,�AܚTْȽ��Vb̙lJr�j&��ʀ�:3�l̫EK�r�&��v��f�K��|��eV� �_0�7����G�ke��>�,����@��o̯ʕ�����^/؄�"6���]��_��
[/ǋ&���.�9�{n��B��Vs��V�C 0Gf���1y��Q�3��?�Ot`�ۧAk`�y�Ev	���~���U���3SuD�Q���z�?J��؎� <�xc��rr0�`��/7pZ��U,��K�����=}�L�E�/vM��=�yɽ+�����h��۾�0?��j�ښ�.4��~J4F�2ŤP)��(���4����G޹��!��e���Uj�,Bm��������TH�~�:��ytT(l� ���hn���ɞ%�
��_X ����*���n?����Nl�7� ������6���E��J����2Bo�;�:@n��K�H�Wa���K~�����Y�N��1��.΄�#��9��\�����a�i�#5Ӟ5�&�LqHKM�k�+��g7_����Z�aZ�^K�@])�(B"�iFN��ȯZh����������o�؅�v����[�2����w4g�mRE���U)���z�4~R�n\ccrc��0�� adHh'r	�N�1P�)]�$ K�af�y=c���ߥA��s�\���_�c�Q'B��z;��5VpŴ�M���Df�O��_}u�v#ڵ�'��m���fP����*E �~�I�jNi��m��T�0^Xw�U۵K.ע��L5j��G3$2�W��hŠ�Y[�4�/,K�ą��_sT�v��JmB$���y}J����C�
Q��yd��1������0��V�0g�*:7�v���K�C1⍛b��N&��6q��{�6[����j�Y!��~B�o�h�v�KU�8�j�0�Q(��t��rϙ΀���+g�Y�=�;�>\_�� ��D�v��2@��J�'����/�x��
'��Z�Jo�]�Q��A<C7�hQDY+�(d�v�t�"�bR�7W�t`be���$��H��Y�;It(��(��K��$���o���\u���Hܴ��1�w��DX�k� �~���:�7���l���9�m]��Y��*\���e^�V!?��,�&��eh��]w�����MK�����Q�j�aN�֝�����^-S�k̢::���QY�5�I�m�����OK�a�;�ZpG�K̏
�7�j�ۉi�ۅ�)�c(�b ����z3	�8%���OgC(�ҫ��-^�8q��'$�2��_	'E���,��7Z�BJ��p�?�o)Z�t1h�����\���)rAq�����ʙX:	�ۅ��F
i\{�1�o�J�ӫ�)�����F�ş�i+,OB�E�{tm��v��m���u�@^���|L��`�dM^D�r[MN�t=8ȸc07���}�4V%{��#���1�z���/`&�V{�Y+�Vy�F7hR���w<͖�yB?�۠n�����U-�@������ >�鄎�L����g��q/(\+%	?]�uQ�o��]�J�B\<�I^�}{h&_�)�dl�J�2q�U���b^`� �C&e�	��� �"��̣����5�#�#�����;��_�X��x�svz���6"k\F;!�E�R�s�m&�<��Q0SU����q��T(3��2��3w#�J�8�z�o;�����Ks��k��掔|>
H�P�T�1����q[aw����G�0�Cy/
Ԑk���C 6���3c��(��>�Mh� �,�*%��c)'�5$�d@-0�$�d�4Z�CGZ�aۉz����`CI15#66ng^��$I,�a��~����HXw�?�?+�������-,��:���QsȰ���<� ��4�o��[}p�� 9�$>Jηq���[�O�k�F��H�b@���*g�nq�9*?Yp$:�F��<�L9����ۦ���ʅp���L� %$	�l��FrK��}�"guY�����MvTp1f����=�=�rWϲx)����a�A���<�mY���.�~��yo'�@:��ݣfQ�j�S���>c��n�inywF}md\.�w\$�zؼ��e�,�8��1��&�m�_ ������Ǯ"���ŌvFoV�>�zȏ�j@l��K��dl��y��X�i-�!5�5a0�+Ԙ�{a�(�L�e�dN���Q ����_A圽��6�Q�U{M:#g���"r K$�]�8^�:�Dd��&�����GI�h���^BX�|PAy��=��\���ؘ����\8���u�߱P9l��hk���lej����޹�����]p9K~3c�
7vx�R3��'%R�l�ba83üu��f? �B����_�iu���y�5R�IS'��b/;A�."˻g*\�O
�i�{������DX�V����?9��!H?�iQ�z��ȼ�O�_ˆ�ʦ/����7���ߤ�%�W!�W"����Q�:��?�_���.�l��4��I�˄y�Z�Qq h�Db��w ���n"����?ƌ+f�� j�	�	 �'��_:�c��'�f��%N�����h�Ԗ�S��w�k؈���f�ٳ�C�m�'�GÃ�]�������-J�ߏk<L�0�o%�O���sY_1�<߬`߅�\�@�u�E�Lw�j�؎X�5�fC<i���ܧQ��:Ѯ��{�����ӚG���\�7!�����$��!���yވCx�3O��mo�!�5|�p�U���J��:�G���,^��ݿ��\�{�1�Ύg��9��5�Qǎ��(�l��>�ڍ��-T���l�#���JH�����̝�#ivU�+t[hJU��+2��X�R��n8��#�ng��\n��^]9��@U�E��V	��O:�����5pnC3�3�.kCZ����rjW{B�mޮ췶�J��aC~+���XQ2
|����DN��<;hV��/����HEE{'ދ�T5õ���m�y,/E��.�q��?86��}����Xw�C֖+UD4�Ӝ�q]L&&(��+5r����������-t��T���v��H�� �sk�!p.�s���!��k�4Mr=�ۀ����DgB��5��C������F>���{���:�I �}wE�D5���8j�`�)�|Ʌ��t_\�6��<t[
�2�#W{�]k8te�L*U�|(�Ivd:׸�C�3,��h�hu�'��5 h�����~YN-5	1�WV�z'��xos#�����{��ր-�FaR
D"Si��ȿ��	�N��[*�* }{�Lk���g-␼��tO�oRj<r�_�g=Kc����"�{˕�I��d����N��|'	@�X�I;݆�pT"�P�eˇH�P��� �2�[2~����U+M�f��������߳z����]�����}2����{;��<�qs���E�#l�p�	��i#��^ၸ�g��W<EG�X�ը����iK8cE�k�Z���?�]LDc����95��N
Fv.j�w .���4�v�4<]��F�%8k>&L\&��v~<mQ9=�*Lc��n
�c%�"��?�E�V�	J��|=���h6�)����_R�3(��d��WB!�%q���nU-
�%yR�3p�1�*,upwr��n,�˘2���r!�����+���A�FԲ���wm��Ҍ�#��Q��0)�t���fR��ĳ"��)�B����e2��n��ߑFI)�n�s��vQ�a�n�mB�.!6e�c�%d�SZ����a�w=��үw�H����P�	<yN��:�Ǯ���F��d>�B���6�/����OįcMݴ��'m.-�ߢOv7���e8*�_�,=%&y��=O���o3�qY����]�oS�bD(��ßnj�:�eI��B���mk���α��c�o!�w�dwt~.H jcÅ^F�M�Ij�FN���@�'�w8�ё��p'-,�ޙ�^�!�O�K"��m����ǥ��3�(���N�X�~<t:���K��L��<H8e�|�����<.t[�el����O�����s�~�]?�(����+I�,w�-ᨲN��~�e��e�R��<1�ayne>��YX���"F�8�PEc�����d�	,������z~o]gą��pC��fW�邲�tǾ�!р�m��w��׉�[��5�b��ph�����v�4K�i!������N�f;6���&�`��.k@nK�c7���?��@Ø�^�񂤾,T5���-�Ͻ� f�[L�r}�)�e޾*�%��ї�������5 ꄽ#�gͲ�$d��2z����z=�]�w�@;.�e�܀:��`���P�z-P��V��ղ��� �Ekv>Ԕ6�;�.����A��>� ��0^"Ğ���j��#���Ǧo�"��40
�J�a�����t�%��yX���2a��Fsa�b��JBn��R�M�� #�h����r��Y?���ӦJ�&Zuы�mP�w�^��m)'O������0c�@]�kX�V���Bub�S
�<���a�s��H��D]$~���SYc�jՉ����sDb�bsF�D�F�g#���`��ʃ������AP^~g_Z�_�cu����ft��EL@u�F���
�-���y�+����Ⱦ����]�?@�|�Oxf�
�-�:C�J�OF�EU�lo�I��$�	�M!�+�$�z��db2Dj�_����w*KNů��>xۏKV��-V�Is_Zװ�2�<�x5�z�+����z���d�!���f5���M��N��a/>�E7�[crT_R��2�+�)c=A�E �H�E���ߔ2P�O,�K>Ǖ��\�[�Ê�+Is�6f:S� �M����]��C_⌀^��m~h��v�;
�C�G~�G��)AA���@����ˣ-�+�Bd�Mҕ$�Z�#���ƿ���k�En���$�XȰoz� Y{�!��6#�T�W����J,��������mwdl'gW�|�CI;g����3X���3ʾ��;D�KX������9�ס8�<�[�kSH�3��Ƣv���e��� �'U���x�!)�	���2���C�ߊ[�.w��&�N�\���8���?�?�A�dw�b:���̜$KHgY*�����%GI*�9�)��5�/����b�ŞP�I#ؒ�L+�n@���yk)w/��4�蟌%nJ�&=T�%����B�Y���;~�&�t�"��Jk�;9 ̏���2����{Վ�g�%� ڞg��w���}�#	��d*g��A�7���f<��c��`�"���z�Xo�HǸ 5����y�#�1�ߋ�ص�%QRD|�9�	쪡���Lk��gs���4Z��V VR���2��&a��c��h<䰙���w_��pͷ#�"��^��uAa�/��ݕ��'�] �����/l&a��O��x�ba���I����i0 T�u|x�`3k-	 ��x����sX��Ԉg����XYЧ!�UVU{۵�),�͹��ҭ�{��Č<,0y�v4�r�����6��+yT�2�����`�C��[ d;.D�w{�m�rmz5�1����ʸc�<:��Y�[{�.���$���H���}:sC��n����!�wU�+��肞��ndA��z�`j G�d�'f�So��1_	]��+��Hv�"@"$�������} Qd��Ǵ`jL���R��J=F���$fiD]��@C�x�[��/ �W�q���Y���,uYpE`CQ����q�IPǞ��P�{_>���*���&�����E��~sݗ���Q����O�/:�#L�/s�#���3�s�g�{fo��tz��rA�r�x�B��I���(A�IM]�m���ϩ�ƈ�'>�]�<���a�2�:�W�l؀���N�fa/�"�z'���[%�Mw��K��֕�ȥz�w��N���u'%�&�:���8`үݴ��<~\(��9���Ж|�B3��n���6�	����u0����њx���%�o�ul��k��%�����R̃pN'5?srR����Y4�#>dʂ�.l�X\�9����Lvi)Ü����)�Q�%���g�4���r��%��G�#�Y�:O�_)G�,�y�,�6f�z*�3T�:�ՠ�Ǻf��b(er�l�o�lѩT#��L�h��0.�,�a��م�����cp♌�R;l��j�j.w��������K�h���*�]�	\)�W�z�����r�
w��d_�����k^ڭ	�O���Équ>�|æ1���j��pXJ�u��I��qG�S�u%�����u�5y�!ٷ���ZЇ�I%��	��V�e�����4��	�����2*���4�y�_"�feO�xԙ�@/��|n��(���Yش~��jAϊ���9�!�,�Z��:��'xD�iS��:��RoF �p-���7-���XGÇ9�Ù~O)B�Ct��g$�����'���h��)a����[Y˦���T�KqY7"f3.ӈ �8x���K�b�`J \��y�(-EC��st��/�t�aM8�X)/�E��u�
b@��,K�^������ [��G��`� ��Ī�oA�:���R~��̷�ۣh�X�Վ%�=�$���oa���7��7vl��ҡJ�����h&k�hsҊx�<��n�����A O�~���`��J��=�bd"!�J�vn\5��^"��~!�w+�#��V&�$�!����.��ÅFq���co�A��"��>H\r��O�y"X�W7݉Щ)E�wi[��tQ�z��N�4�a*�1�>L�c&���@����k̗)jLb��?�:��;���%k�<qKZw�q�,����4���~n2���&����?����T�@M���xtj ��DL���J�z`z�4���L�W�dNJ��0p�\RO��Q~�X
�ޮ����K�S!G�`���].�ZN;(@�Z���CoqL��T�aĚ���g���oq��{+��������+�6�Ubgz�o�(z;��q@B�x�,�P8���IN8�I�yn��g�WT�+���<�۞�����r����v�m�	�ˑ��%Cxf�sVÒ�{m�:U0�;�k�$w iG�.]�Z�����;���0�����y-�7�c4s񇘺�O:����Q�%*> ā'�U���k���M�h��[`��3<��"g"�=��V�D���*ɷ&���0ITK3��G��߳OS�>ko�:�*��B���v^�L�u�Gy3�Z�b����,;!�Z�T �Q|{< ���q��fIt�5ڃD�{plJ�f�,W�Qc��@:t�Q����O���m��S�<Ej�@����m��c��'ԙ��"��V� �5[�Ѿ]��&���4h�*4�j��0z��{T:�Ѝ}dhvN٬�RR/
̈�p���%W ��5�;�E��V�q�w%%R��B���w���r:��4-�B"��뾤B.'����
�:��eB��w����	d]�(Hg���~�==�f�1����%qR�˼�D�a������!�*u�*%�ڏoq���n�i{m���AFu*���XzI���4�fc�����r4�ACf��5x���$� �;1Z�dr�X�������@��Z�����6��������ռ����{R�o!�w�笽=V@�0�!<�ܳ���{������hW�b�nB��'��`Fd`�2u��r	~ o2����ڒh�E�b
�_�\A�]�e�80��-���}��5�g)x��;���6����� I��Ti�����-�9�_/קD��C�{xŲ���1=J��*��N\��'q�V�|�U�I���b2=��G���?`�L��f0����9�;��(lm6�J�y���/f%�:I{���F���e���z'-S��*}z�n�������1���q�O������Yվ�^~d*��ո��P ���0���)�3/���/ O��N뫟i��2ɞVYL�0ݾ�+@�e��8v�%��֌-�rD;���Ow��:���.w��I'�s�ZN�T����O,�]J)#}p *�X]w��up��T<�ˍ��A�f��)'�BX~2&4X̀W�?�������;�`�F��%R��MI=�u�b?��~:/*|�Cf�]f���V�;
��j���bWV��YįF��\-�?��ZA5��ݛ�o�5!��'���:{�m?c{������0aß�u�4N�0��I��φ�<�^O�VC9Ll)G;|T��~����-z�"�V���Yk^BM��g��A����J�h�����q���VV��h�.^���&�I��^L��@���|�����Kb���q��R1��-�>U���,E�ꗨ�I�E;i䨡U�xjc��®E������ �A�j�d�R�L�h�O�2)��`j�V��<Ց�^L�LAm�Ԅ����H�����9[���5'Ƨ�͌�F���2���~�ka�p�囡{�*���E�w�����A!��?�\���6Vq�b�f?lK�H�)��6��"�{U�����3*pE�QLZ�o�?�5e{*q���Lh͆d���u��\�-�%&P�#B1I�ͭ}���8@��pP�օ��y���%$jZ.]S{8R}�˾��q�hjj_��J�=,����4���@�f�Dp����;LG^��U]����~ћ%�?�(�	x	ߥ��˺^H�O����2��T�!Q�m7�9Y����ҌM�u%Z)@7�a�Z�H>Oݘ dO}�.�ls���|WwYۍ$8b��ż�u� R���{��D�G��J���缳�#qE5i1�!�G�W��sO ���H⊃�v��; 
�:Oq�����':"[�(?�R��h�{�K"��7Ӿ�,e�8�=��i��>d�������)|0?��[xI	�2�ُrw��Ii�|��MT��{�뒯�ARL��^/N�b֘�X˅{*��L�z��r���:5��\f���&��H��Fф V�~�<Qk�~��癗0b �YR���� ��x�}[��I���1Ҟ��k%J t�?]`;��X8O���4�[�-�f�2s��.��`�B��FO��ن+3�झ˾�<�w��V��zU4x��~�kq�aW�?�) ŘVO�>��#e��M7�<v����?峘쭰�Y��`E��Y4�7��݇�ׁ<+��R��R�F���Cl�p�'��q*4?���%n��-N;V�YdӪ(d;���㄀;�r��=�����
4�M�BK��p>~6;�j���N��/��$��G�;�G���hz�B?���#�Eqe�v���V<�-	٧EՂ-\̲=�E1_h�+�S��1tB��֧��|ݴ���n��/&G���­�`sϘ�gԲWX�O�V4KbN�34����7>-����7L���ٜ�@i\@�T'<�`bP��z���Nk}\I��h�RQP,�>���]Q+ gV!^�w��EH��#Yu���`�D�/��qæ$\R-�i��,N4q�E}�[4�0JC4��r<�Th��R��/���f�ګi(@1$�ng�D��^����Z`M�f��?�&�������]���|��	���t�b��� ,�[��ϑ�9pSKb���&�U�A*�;�z:1�����֎`�%D�,����-�����e8��e>������6���b������+��^�c����U�T�,,Ր��a�k�5�3u������]� ��xE�m��3���~���Ч�y��܀R�;yjjG��i��F�v��_��mC���qD�ȝ��l�6���Q�*G$�>`<�
.�.��]T�+^a"k&`��Z���с��S��'��*-��dn#�+	�6*�pD�I7u�r�P����Z��ϲ����w���l%��7�oh�Ż�B�����b!:+(�
P�Kj9j�+�	N�@��������Ҙ���J����zQ���(�y_5`}.�8�*@���dz���X /M,5!���(�{�s����W%k�es�d;�@L������l�^�$o��&�/ͺp E���x?+���ND�n���˝)�*VӞrj�8�Y<�
��lC��}� �߲5���}9�Pf��*'��~,vL�o63lab'k�k���3�:���³R���Ul�J�<�[��yɳ�s��U���獊�T���U6��@1{=T!������#�ڒ��'d� ���c%uS�tӦW�Gj�v��d&�v�_�b#&"��e�sH@�e�L�-D o���L����hV�b�m�-��/|7Oe�m	B��R�ƙ�}�w���(�����w�Mt�����?|%���֗~i�&*�az��mRVj��F>�{_s�C"v 1�.��b�zD�k��I��N��J��1ꎉ��v+Ӻ��8�c����t`����-�\��I5&��X�HlR�%!Mb[��g�@�,�*�]"���*@�\�3��VM;\�~$��G9|fe
b�>���Ƣp��������i�x�^��#Q���50�|����V�3�-[>#4� _�xs:^�P�e$<8��U��%l��DE�8Z/�h�=&]�nzz����D�^�Υ	"\Scl�7��+��讉[�V>�:Ơ�F���Cq�_��ǎ�-���=�������M����C��͒I��A˼��.&�5�����̅�B�Y&y��t�O�tKz�����a	���+z���}g�A�md.�H-��5Ql,uQ�j�V�/����Ms��y�ħUul!H��s/K��kC?�z1���vlWu��<�������go��/�Z�צ�R��IH҂:c�1���2� ��-��mr��F�6ZG�*�?�����[�E&��J������31]������ׂ=�"�G�E'y!X|�����	��asA� 	��޵���?�l�Y�n�˪��D���S�]��Ǻ�h�Gr����h m��5�;#�7$e��e/�>�bŭӎ1D-���cSO��)|�Z��i���3��G�N0����7�j;�	fe�O�+���ｃ�л�f3=�	X$�	��E�8��k>��@��7H~�M��8mR����;v�~�J:A���WV���.��ɼ�;}�����ɧ+K�:<����X�U2]S��~��<��T�Z�e�x�u��k|�^s�`s�BX�����-&l�߿-t�HÀ�RjԈ�3�Q��9���$��V�`���5i�g���o��A[[t�b�ѡCi���l�0{F#�5�;S�?�	^��<:��.��F(���q"��U1���1�~-�?%MS�i�z.�����F��B�r�Z^X�6z�)�Έ	q<��_�Q�Tc/S�9��N����^��ҹ�&��)�	e;�T��>�~�2h�H�aiտ<$S���0P�As�C]��3̣H��%�1���XU&0[�r����m��P��+S��р�ab�h�6U ��UF� ��i�q�SK�C8�kyW~���k5�j��#��� ��
��}Z�n�2���&���W���[���Z�s���=d��u&��^gCM�#�v�����zL��^W��3R=�zR�Һ� �cgv����l ?���T��S�jw�4�_��y�Ar2���
�"�F̵����L��{4�s��1=�Y��5����._F��R�>�n�����YV\��M��HUz/G��ʃ�;�q��H��]w(rf��x4�ռ7�9s� p�t���c".�x��q�hͩ�|�W�@Јžh	d?��gSv�Ǜ`|U�_C�;`/ZO����x���Zm������U8:��Z��C��1�i�_c0����8��6�4��lť�)wI@#�~3wVkQ,>��H��&��.�T�K���M�޷8�)s)��ΩB��?X�٦���J 4;��v��=/1�X犨dW{��?=�OXz�w�{���|+��L8d[�W�?m�"�Hŷ���y8��*�׏�~&�rv��Gs�VA��ݙ��S�i T���IwA�����;@E?+ND�l�䙐�!j!?	4�������٬�qp�]c���v�i���/?�=K7��[vU\���m���s�i*��ciذ��1TEn�.u��U��-���9}g��u_�D �V��}�Մ��OxO�|�]��u� 0��Pk�-�p
b@:F�b|���x������w�K�R�Z�����3���Uu�#��:P��Gx����F	��S�)�Q��<�R*T�*\%q�"�B��[�X|Я��7�^$iI�;Pv�S������_�?��᛫�f�>?�o��G7�
�� ��@E0��ˀ��%+=�V]��Ƞ��Ő_��a�)�=�<q�	@<g���J��/C�m򬙼*���v5��5��/��B7.4�e�6�\Ŧ���[����֕�(�坤���tԕ. ������� ߶��b<)�ma'p�]m����1�~��]9��6S��@���'�Ó�5 P#���-'�ě�՞�ێ��$3�!��$�*�+��Fua��0��l��fh�"�X8�*���.�<j�x�I-�Qt�c�G)��痍.��z���Q�d�/mѺkd��Ȼ���'J���c�e��=���87��F��x�~0��E'>��}��+��#�Sk��e��J�4�Da�$6-^��.���r²6n���_���RC���h�/���*�,����q2:�[`W��#|�O���oݴ�ƌ�"(�xB+,ģBT�}��l\���#�KJ*� 8Y�sg˹$�-tuc;�o��2�/���r��W�B��w/g�pζ�IC��'u%t�2OR������k/�p����E�y���X1�,�8Zi7�]�Lf�U�I�彼���~Π��Ts�/��^rQ,�i^W��5H�o�Ics"0(��ab>��R3�Y�������4B��C>����Y�* ����'-+�s7��G��A>�H6kR-�ܸi�ؽ��ϳ5#n�)u�����%'�Yl�l���Q��!�]�^$��X����W��°ylÏ�+�2��	_U�s~P�[b�ոv\���**��!�GqD@�6�L�2"���.j��v�,�(�+-$ t�����᳠y��YG�l�����
�m����J����l���|�6�.A���&�t���u8�P�^��Fb	�"���re@Ėx嵐qI��e}�:�@�ŝV6�y{;jFC����E�G�?m��M��{�oy��s2����������,U����3�pY���M���~�@#�����^Y��M6�n���� ��Y�(�|�����`�?�6�7)�U�) �m�fȎ���`gݑ���@�E����`ٻ�9�2�!���d��	(r����F�(A^�Y>$���B���ż�r��)��/ؿ�q9#o�$��88���Vmsmѱ�F����ϴ1�n��=�$v"���d�us���=�E �{AI����|����� �73]�m0b���.m"Y$�e^�����p�ȱ��������I9�>b����;1R����)<���z�/&G�_��ڄ�zs��b�#gh�#���y��b�A,�^�?&��-sn�V/*�""43X��\��$g�v*�v��q���&tM�ݫ�@(ͯvR"7˻�R�f�"�A�*�#GPX5^�+��0�o�s�����Sa�C=�ߡ{#(��`=8k=���/i�6����������
%�!d�h���� 8d�����)�~��
D�i�&5	�'Ur�!�*�a��@��[S�˲�"�M�◛�p��xc�����k�^�5���������o:�>��n��NoI�NB^�iu�#w�Ӧ����K�
�׺UgL�M�r�~DL�!5cb�"���M�gu�0$#��S?��'����P��%�RM����,=K�uo��\kgߪզ��$���~rH%�O}���<�ß�����*GR�+�VZP$�輾x~�zf��N�<FW:�?����3M�'��;I��P�0��t�`�M��P;�̒��#Їƽ|8�W�W���
��9�d�֊���x����Gb�De�R��lK�e�_F[���S�m	�E1«��V�m��û��-8�ÈL���Y�R�c�D�����2rBN�"zc�yQ���
�a�M�S�(,�%-�w�]Ƃ�u6�d��U�]�$�-Cr]���r��x.4���ϔУ��EE*rb�������{D�E�W2�K4�oi����1��7�V�x���=�!L@yd�� i��:Uq�5G܄F���L�(k3����xp�G�xB���Y.��g��
���	gTȣh	9�k}��y�IJ��Q����^��i���('5�p���i��h��!B��A�g]"X8���E��&�kc\2�ķb:?9s4���a]&.�_��m�H#�Ńz��8���W4��1�ƀR>I�B��==�!Ң9�\��Ba��Y>L>H�X�ZF'"�<g�,X�ɔ��T}j}����虉-�n��xs�ؕ�@�f��l�-��(� \�>hIB\'S��U�0�R��� t�_3��5%�+�,�kRZ� ���-�9�O2�4���Y�1t�C�#»�U�́�ٳ%����W�a���'�1��m��$�%nH��xS�P�nHr�2�殞O��jg�Ly�S|��5-�y2f�~#%�|��-���gh��R�����	�N˵<�2�������"�tg��R�) BfL �~�K�VL����vЈ=��F�?��9˦��Mm���'��=�a9bt�Lm�G��z�0_�M 	H{N���JN���d��c\�q�Y[����3���1�F����`.������s����>��Q���[�,B��ChL�l���d|�T�[��^�,0��������u
����k�0o:i����ۇ.$���%!N̒Y��Df{-��� �5�6-z��#�@�q��2��);XQ�z,�C�P7�Cs�-Ap��hӱ�)*�$��cl���PC�k8:����f����	���3=����PG���//����åQ�blS�����v�/��L�WӥEYk�C5��fMqe���[O7�P�1�ӓ}S�f�˅E�P�x%��*��	 d���~��������KI�[��T7��ġ��� й��E����Wy� V���>s=�/��|g+k�c���=ګ��,���1�\A�0��[��L8\��4
���X��O�re� ���H&T��M*]
�+R��2?�!�=1�o��'��)��[���}X�^ =�G5sg|�M��oǏ�c���^r�b�Ř/�{%zљ:ň��N>ie(Qm�M���M�_�+y�Ň�3$"��WT�Z*\z4�j��kW����#�H<3�^�:ɾ�/�Y�tQ.*�������T��~���u�ԇA�{R�*������M!�:)߄��M�t#C�X�U#E���:(Z���[a����v����դ���	�Z��� �rn�5G�o�U�����;��mh�hXr�#Ҕ��ȋ�g�'k�C�)>��L�\��l�ﳑ�M�i6+�	�3��W]��.>< ���U��1��;R�� 5�S��� �TDG^��o_f@��M�m��m��ͬ@�cf���p��q�`|)�$\���)������i�"���oXg�;%�}i&�n<h������Ru@~�5�I�JGkK*l��T�n_�m�nR<|dp��E�ؗo���jͥ�K={g�~�@(�ꞃ���9 k�	m��{�^f��=��?��3�F:�g4ϸ �jv<�Z�� ��
�)�F�
����d���{�������o���3C�C�#�V�xݫ����u�b8֯7	��g���TZ_қ���$)�\6��rD��D� ������iQ�\�:�g���
�c<���"�sS�!9]:Ϩm�{JH2[��m�8�ٯ���[<-)�m��`�� �1�̗" �P�§p,Z�k@be?��J=�p��-�KHu7l�h�@�J���hݓ��?y�i��a�9�����X(���	��uGbTt�ԍ�
�	}�	q�k��^�,.�	��i�vt��A����z�&�x��>������$�Zb�@~}+�q.�f��U���s�2ͮ����0 �m�R����/}�4�:m85�*-����
1��M�70��\w-f��j�z=Sd	�7z�cH���N��w|dn�E�݀%M��R^������X�N����O}�K�j������_;����$��~�j�걬�t�w������T
��Z����߾�ӛ�j�٤��nn�7��*��KBn�Y�9 ��9�����~�P��Q��u�r�@�{K �?��u=��l7�K�9��7��V�	���`�g\�s�h�����/����jK�U}�cK����.��H��$�N��œZ>srBR��������\\9�(�כB�o�Ͳ tK�F-d;�9�����v���T��$%�l'�|�ɥV�y0.�sK��e��\Z"�K-~��05�������T��/�0�%�O��\��v�ޑ�8L|vF�䋹%>�C-�_���o�Q(�[M���2/�E��2�'9��F���E~]n��2�?�>.����Ŝ�U"&�dcw�M��'.��@�E֊(}t]N��P��:����*�z�������܍vҍĠ�dX�N,
g�ExL�P:4#$�#sI��iO�3&���0�9+O*�}�\���xMDo��W�Ba*+�;��Za�i)����~u������z3��$�	|#��-<V���k'��3x�_��c�Q/�h]���pt���ȕ�S�����c9�Җ�ʯ��|{t����>ٟ�ë&�x{{5�,�����X��� ʹ�>5Gx��%�n�_ �=���]�Z�*S�" &�����>&ղ^D"Y�ib�g�����D��p�O��tt�d�U4J�f�LI4ُ?�-yy�.{��h�f��cZ����k�����ȉ�'��w��g�M"�_R��vI���0~D<3	���pGxP�2VU�EWdG(�8ꓝ��bBۚ�ܗ(�!�$ �/��F�E�޲�dq?�o�h��9�g��>b\K����J�%;j�z� ���*��[_�5�\�I�̹�mXA)&���)�R&�u3�U����\Ck�P����K�
�zs�b.���8B��"��.����:�!9`�7G�7-
#w�<������N��D���������=w�<�J����k��T~�b��%�ĈI��'w3��uߛ%0A��N�43r�9�j�7�ؕ���`x��QU.qh;X�ψ��&�6�Qj�H��>�?~���J�:@�\j�()֨%�� `[t �>�.�g��+���<k*�1��:�i���)����z����r�|�/ͤ�
YvB��7���[kt,lJ9�!�99��J{3���44��9.�@X��Q���՜�c��%�P���CQF ��28��B�ў�^�e.W
�0#��p=#ښ�r�:m��s�ARU,  �]he0<L{�V�B������ob��\��&/�{�3�����k$��#HMR���e����f@��2�雙Jg�h���BЈ���W�\��7�>��5�Du �}>z�gjڻ�!�]��W)�<%N�i6�ۛ��ݥ�+�ɂ6�p�H����vĈD�9���5�w)�f!�?]�W!��Ƕ-�,�>v����B�(��gI����Ee)�3�UD\,�h^��q�R�&����;`K�3�7�
6!eZj�"���������P��J��2:����Lc�{��<'[u(���XT��c��~�;^�!v?v�%��kͲpXR���Z��襋r�-b�ȑ+�A�'Z�#���Xh M%{����P�z�+�c��$# ��w��c���6���b����h��`�ʆ��l��ycoh�Șp#Z԰keucg��"¦"�uEy�/2�����6�@����2H'`��S�r����>f�l�f�M�{FՉˏ��	|X�`;�b0s��@��N���[Z;�û&�϶�Ծ�K�	�k�r09p�����e�%�l47� �74�u ���d"�J�	ކ�'�����: }#�Fr����&����i9Μ�J�p�A�r� �~
�;H��Û������pdH�x�N�z]��!| \L���� %q��
4K��{~]�H�L��hb/)CC$��y����:�j�ʟ9���Y)��t6z��c	�@���A�����e� ���9�D��J&��4�$wh$��t��y3�!+Ĝ������\Ь�M��Y��#܂�Pxj��K//�Ww��?�LB�dF�U��u ��z�T
�TQbe���90�p�ߺ׋��f�$C ��i��Vl1�'IA����͊���n�cx�V�p��ߖJ�s��d�=Tý�3|P��c�K�`/B
fdj7G���I��V��5�'&����ڽ<���_��e�O�X��,9ɿlӋ�I���j�xpP�Kϼ|�R̓P�ߴ�
2�¿$���+��Di�()�6�XiL�e��i�ca�G��>�p�LT,j�w���5h�'�5n�)Ѭ�0GD .������C�)hh��$�7I�Vs���Yp�p߫�u�A��K#��s��:,��:hϗ���i���q�����������1r�v�:�\"�G�"q�B��r﮸_�'sa�Q4Ӣ(>r=�t��-�w$xSS��c�+�埄��#�;@C�gҦ剴5>����b�������(�9��OZ����U�8�8\y�W2�ߢ����ڝ���mG�:u,/��_[ Q�|KLV'�0+�}�~�T�=s�B;��s"F��Jp���bXP|����p��ƫ�k0����1�f	["dq�z�hr	{~�����P���ۘ��ѡ.�`���1�4�| �ݖ��יT���;x��e�Q��{��.��!����^h������%!^�|�C���,�E	.�<b����$aa1Av�0d9���E�,�b�\5!vk}V�����'U���)����ii�T&���`�)�\$�W�j�ח�:�.�6v��ƞ
�Jy���J��ٖ ������ۡ�:<rjr�C�F�/�S�ԕ��g挿��o�Qd��? �^y)\k��_vtN�hݖԱ�K̎m.!����3����= ]���ui�׀�x  R����6�g��^��%�^�<�H!3��9#��^���Z��՗�[|ұ�c�a�����!LO� ρ� �
dUh��-B!d��A�3�\��]2}g}�r"�Ι;N�q]ۮQ6na����0���Y*��p�����ԗ�m� P!��ZI��0���-Qm�1I�m�VV^���A�����$����&����7���/9�t�Yr����Lr�D��T�oaj1u��u�msr�I���3�ki�6������8 � ���C���: ����H�bG�ozE�&"���v_�Qf��3�r#��l��(��4�3	e��ѣ/���{�3���S��ׂ�;�\*�"N}u�[<핚��Y�n_'���'�/���f:ʦ0�o2����~!���;�o,���'�6"SdP�>ҭ>��m�B�s�(ؚ�?����MKj�^��Pi�k�U�������)5�cv�ƍ�(|}N�+>Ąnﴃ*�r��UU�=����L��R��Ci������[ݽ�1��5�b��$�D���U��C���?i����j�逴N��A�X�<a�0�C�5�J���d.�1nO��{���G��<� rd���ɓ`�Δ�NlS�-�.Δ��/ǔw�+���Xb�>Þ.����!��(�c-�6%��C�*��f���+�ǡ���[%A|�G��+�u��������ν�%���qs�	5s��^"[��+du��v��V�J��-k�ec���K�	I��[��6�캍h4��C�v9}��a^]5_�F�]d�sG�l�+.��*�ORz�0i����b����f�UW�G�.�'(�/}1���6���L�x�OvS� WwLjt�ƧFW�O��y���w�*��3�C�3��C�(m��E�v𜊸�:}P@_sY�xt�k-�g,��m�ߎ��։�<Ч~'���~Mg��s���BpF�}�j�&q�u�&l|�'(g��WEL(��r�j�:�D����n��Z�G}%�wA�ٷ�NZ&\��8��EH�T ר�h�+��:xƷ_	��t3T�Ύ"�6l�z��T���BK���y�3tt�`W
�"��o F���pو9�}�����>v~��U%�Z�?�]�uH��r����'7�_	3�����I;�Ć��]pB��Лٞ�SB�a B��J9�ޅ�`�w�A:�ѝ�AѠ�zڝ��������2�f�\�����v`c^���lZͯ�^x���n�*:�@�h9��YBK�&��ԍ���z���F7VcY����@�?��hq���Xb6�9i}l�Ӧ�,�a��H+��ZFl�w�z�]����_�����d��1�PH�(�}#���h��Q>ei�I!R�����1l�W���7�غ�M�f�jʟEr�XHA���7��@.|��[*����U��h��^�������,cJX�� �� �$Zt��<{4y�ѱ��KB���r���4�� o��o� |p4�lj��/����A���m�z�`�_���U�{M�c���:��+V�a��sH�7�s-6������	�#\�&�]$�"�tl����%�k����-��7/����u{�2w�V_esP��;{�S�'Sb��?.܃x~��� �������6V�w#���Z��l�/���*Y�A���GgI�n)�˴AH$>�L��s�T�����I����C�y{�N�)�r��O,�����KGA�A]���@�<�8�pNz틫��a�����6��ۑ?u8m�P"�K.�,�sq��_ߗ�퉧6}(�sb�b�ٴq�$X*JK�M����a����o�sd�l5$q#��._��ܵ�?�	-�w흍��N;qj�F�-�T�$�W�H�c���"�=�u��3��Z��֓�P��aI��"�y�n��t�eo�9\M� �pΉ���}��JR]Z�3	��ä�Q��`%��3rCgT�Se�ǗB/����^��Hs��]̳6bl/��8@��;�
ф��R*V���}i��C[��p(�&*�C;���(���YP��q��:�!ӹ�܋��ܻ�9˱���ġwOa�d<�k�h�XܒҮj������}>_'��� ��^�;�3+cP�5i>b��O����ؕZv���0"\�ݮ�R��~4�xǆ!ɭC=4��J��PE\�nہh�l�개ҫ~q��=��3u
�Aj�q�#��>l=JG[��o0��D�9��Z��'H��+ô�����\vҞ��jt��2+�s�ƪ�'Wq$Q&�'f����wv7�ƅ��z�gd1A���Kot&��n=�m^bJ. ����vhG��6V�ۚ��;��&�Et�# E�d]�źg����"-�{�m�Y�J�6�g%�T'�`�Mk�!R�\��E7Z��i:�jB0(p�j�HL/����,q?�ѿTRT�V�mVC+-�8ud���he�<�5r�$5.B_����k�9������~~�.N��k ���뤓�oF�5�����2]�ظ��Oq�b�u�"kY۩���'X hX��`7ej��W�K��БЯ�.7���Y��pteД��у�T���E��RZ�\�݊��8��]w�^JvS�������������$�\�m;�+�~��X��is��%`�Xa5Zf��*G��[f6�b��xa�њ�{�$^�L���#�>���'��%�`�Ժ]`
͠���x��'�^�T��1f�������
��3|�;�#P��
'���y��<&�^��ej���"�[�K.��~m?��ă�[�}����k${��wnr�\����������aPW���2l7�y7:�ԍ2JPhn��lb��bv�|Uv�m�tT���`b,����h�J����P�S:1�(����Y��V��B� �����P�n,�+F9[�s�;�h_���?�Єҝ�
����,=�6�s"��1+�uKu�oyU�M�f���s\N#�sܜ�r»�m�<�u��ioі$�ɯ�g�@��ۍ܄W�?��)��s�U�,�K�(�[�m3�hk�B�\k��:��P�JH�&{.L�P;�J��v�`�Q��?y͓Z��V�r9A����h1:J���ڂT�"���{�-�:RGjq'hk����r�����f�r��d���}��)���L�\�%�w_�A�@����,E%�	���6��~��N���p���/�UT92��۲�r� ��5�my ����Q��FH�� �t��SC{��� ��&��<�"}�z����,v�}�\�d����qU"�#�EK��t1H���/*ȕ�4� ��+I�Mأ���0N��Vui1�{�F_�F[�7�y��K�1��\���h���1�������.Z�y*#=!��Q�����:˱�� �S�\,��,9�D�U�Ɲa'�ie�%�h��l�뱞�v�b�=L�F?Q�]��__�R��	fڐ�]+�ax܄  \g��K=���J;���_�!X�4KD�h#���7��Df"�J>C�4��[�]������ꁐ�_[�v�6�6�s����ON�@5�/�.E�x�}��U��LR�[{L�.�!�$C��ީ���C�ת;}gʪɻ�ӟ!(w�P���'���<DB��o������6R���t�,ޚZ� p0�}�Xh���TI@�:{��^�&�1.~P�n�5�aa��Θ�6&)0fo������9m�&$�j�c�U��I4��x��|�b�����1㤦H�t�-b¬6�!20�?�����ˍQ�Ec&�9V,�?]EFJ[�I���ұ�}l]3�@Pk	�h� ;8��g���ܾ��{$X����VB�SpQ�2����C�)����R7�O��@�û�����[qH
Z�&�Ԩ!L��}w�8u�p�����Q�} WP��f���]�!��Kq�v瞎�p����z�`;&
Q2pw��{��M>�>�ʫ�������IO�@�P� 0��L�2���-�N��BZ�@�?q���
P�5����(�Cˁ���H�	Wc*�Y��M����@��!Fv��d-[�/DXH�QS�}φ��� ÂS����g0��F=���P.N��<����`�#Ps �a�����(�T�٘\�S�&�G��s��<П8��^}rAS��0q�
!�;9�r\�&|Ry�8S4���r js�x�W�q�2�%�:����qQ�I��5�(&�stϸ��o�:Ĉ�T�A�l����z��=��p�j,�-�05n/B�S��UEm���,i�ۘu�K2�����4
���g���#�%K��P-o�o���}h⋣W�1
׉�,�yW�thD#���`�C�{���P�r�;e����Fv�?
ٕ{�*��s�6�VZ2�;!�*#3��H�O����Y�@�+Fɩ��:|֮�_']S�	(b�!�?~{��c�)W��iE3imP��}'+k�vloIc��_5F���iM�F{�隸��o����o��$�5��9h�^�_�USEx!Akd�����+м��3^ƋÁ2�HO4��U(f�L%^���3A��*;�`�h�#��O����/2�?F>ǲ��|=�6�6H��cY�C�����0�u���0/VC��r��ҚV�7y���k�I��PF�/�/���ש��E�^"��v��
�*� ��W�!�:Ve����e}�ƥ�%��ډ螫�+;� �c�r��	�8��?$o�;����������)q�����g���k�T,Ap~�#���z%>?�K�-'b��+\�Oo&A@���|���)�Z���2�e�a�^�&ډ�9�>s��ݰP���_�qX�*���܅'F՞o���+�������C�Ma��t�'�W<��eHd�ceCo?�����.�6y"�KI�M#z���cD���͍�Z[	���C�XFX���N�%�D�F�>�C����hF*�R8��,�	Xd�_�T�a��+3g^�Lʮ��K}r�t�֯4 �kIO�
Iݪ>��Qeb�g`�<p�uUcג�b�[g�X�ĩ�lC�=�K���C��&/��1�X�R��Vը��������t�0���#h�14/H�
���&OD �M1��B��Py�]HY��i~�5��ަP�y��n]!�\��7�1^���;���b���n�qB��C~��\�0ZB+�фb�F�e��4��~����k�מ{��{��������'3�z�%�q���X��!�;r��)��Q��Q���ȇ_ud��o����8W���v.s.��&�R��.V��lk��s�������[K����O��5�q�h�c�^/��F&H�˺�I��J�!�pC�cc��S��񍘭S��#N��8�����"�T-���7���7(��a���ڻbWI�U1q1��5W������l�f�<�ˆ��QݧP�W=t�#ϵ�D�[6䮷����ܟ ��]!�?���7�O���BwϚ���%��+�D�2��y����}O<;ܜ߰��F��$��Z��9��FC~�>�M�-������.'��8ݦV�jd2�Ko-�{��I:B��2�C8�����LL.�/�t��I��/��!���}�5�vJtoY��o}qCk��O��^3��J����3���rm���9ӕ��E �m�����|{_A�<K��S蕸�Jĭh@ѡ��H�B���w�@�I��'���&�OS�~�d�HfZv[��s6˗��:TC�f�L}с��)�.\Z��uұ��h]D*���k�KأE/n���ms	wG"n0."t�0�N;kl��eY",��=�Y�� ���uw��8H��?�����\ݙs@jBs?����T^�X�㚬��5iNv�Ɍ�eH�����y�25�s��N2����c�7�(�<w��渰�7�?�x��R�-�Q\k��Z�y3�4E܈�T�(@�:%pcқ��� ��l��t���V�\�G(DM0�1�	�4M�G���@��07��wރ�3[��c�(i�R���.M�m-�_+��ȳ�픓�X���`��K��i�0A�rCDU���|^��[�@�ZÑ���Iw[�8  �h��[1v��V${o��v��������̚8��Jw�s�R�3���㸣4Ø�y� �N&[�+���D�E�Ş����ő��K~�����k*c�d��s�+ft�:�~��h
RB��b�����=,���{�о�J�nb`Dڝ\~T��o����y�DV��� #��2�q�wK�����xpa��Y�"�&���^r,��LI���2R�ٖ�$ϓ��1"Ƙ1���/�����w+�+&�.�z��.`=N��ⶾ�e9ܧ.h��Ӊ�T�3��Kg�l1���K(�$4�E)p1�9A��?i�?�f�u�?,�3 �~�`�\;ߕ3t�/�����.��;4�f�~I���3�=�"��M��Du����;>���@��:Q�h�������0 L3r�S����l}�*"��%F`���p��/��ו��=��� 8�������'rL�b�z\��W8-���P�� �
��l�v�M��PZ��ι�D��9�_��G�eL�B�f��yg)}|�(�%#8�"o�i�F��|�9PM��w5c�-�)�����B�j��2o�9�1�¯�����s�z�)�G`L����d)�$���N���)�c�d�sh��K�8�_���������G���{��E�|!�D���0����t<E+ ���<����lK����R˶��U&�{��dܑv�G{�\o�mm��~�g�G�[;t�6��#�����Zu�e!z��٬+�b�N�<��'����\�ÍX&�w���J�=�u�2O=�+.N�M��p_�����41���ia�}29�?���Ҵ*��96�Z�\G���y7�<V��������������͝4p|�r��1��d���S��x�kVQ�gjE�	�[@
��t�9��ݷ��\PX��]�K������P\�.�#%� ��ǋ]C���GH�FDռ�w�4'��m-;�hNal��P��"1�0��䯹�^��Jע� �;6��� 956�s�[�J�79g�,���}���� p�l��D|㶂,�"ZS�cH��3ڈ��**Y�cR[i�����f��UV���a-:c�"�%%�^w���wY�PJ-�b�RׅZLe�\,6����1��c:M����$?����G�[_]ڍ��>�܍E���X�F��2ba�����f�[.r��)0�a�e� ʡZ4�s�V�p߫8������K�`�2$ӱH���aZo��2ݝ���-B4��S��L��Ǥ/�rX��2��;0÷��.�Ч��ZBÐK`'Z�O�h��p���pz�����4�����������_�w�,�/zJ�T�������%�T7L��0�[s��L�eÒ6��V�>�h[�x���펟԰#��\��6.H@!�)n�t����3|E�J3t��g7�[CR�iZ%��f����&���q�F�)�EptRF�����o���x�{1U��@2
s��d�N�y�ߜ4���]�]��d���� w8�K��"���
:�~0γ!Jd�)�?���d�g��%���?N�����4y���s�˫&� ʲuk������ڷ�d�3����7?��jNκ2@R�򈄼�_��3�M�s�%;^���A�z���;I�����C�Ȉ��6Y8�\(�i�s�dJݿ��-��o��+�d6�`s��
������:f;�sj�?����m��DN�,���+��T������N@���<x~̨gP�}��L�g�G7\R.�-}�4�fpK�N�l��\�~ac���0i�j����Y�ͲĆ��q�)��Y�H4>�}�k�aK���0� h�q�"��*��I�s��&q���9 �Lvs7"Եmu�M��v��H�4�/=���$$<�������3����]������ɻ
5��Mz�3%�E�`�H�f �@�[T6P�Z��Nmzɵc$ �
4aSD[���k�����W.ܑP��ûK��i�v�Ns�Oe_�/s�횕��Os<���&�Kk��,�1c;ΡS�xR!��ʂ�u����D�6����4������fG��Ov����ޱ�!���ޕ5�t�r���n[�)�RIؓcr��e{Ȣ����o�_�5PA⨃���2�1y	���V�V�T��6��pW�U�
s���̭qK��4q^�rfg��qI#��bf��dЫ;�\��W;A������r�"SBMI����Ϥ��^������9��M��_Yϋ���ͱ�F,���v�X�a0�\�ˣ,)D�TR����
�W�(�«�4mUb���A��5j������,�$�-��w}�>ވ�JU�
l���{9XI9/��죶+9��>:��!fQ� �:���\��A%&�7S�%��+p
�ckxC?�Y�Qi�����*"��@�'��wc�K�t�;ec�\	����!�ͳ;����9�ܣ�$�d�%!���\�S�t`��7U��"{�c�ܚ�ǿE!�a���<����3�2f�[�&�σ��ܗ1'rbG"\�9 �[�U��=��S�p2ᓁe��2 {J�ns�F��J5^��G�5O�s9��o���9��(5��� =���g�)��(�k5sE��X��?{4�.��˃?��aک��6�V��=���x�E��ዕ�#�$��Y�����bb������� B������.�q���"!�M�=9-�I&Kr6/�j%�i�gP~���������\���p�Y������`�ev�%ӂ�Rg'U*�v �o7��I�Q�?��}:�d溡k��@�7V�7nh��T�����S|~v�Aї!��(���i�ޘx�R�g-�ϐ�nh��]0~X,�'�����>)4�tϥ����wZ�^���F�l��>�6a-x`~|RC
Wa�ť"��t�U��!���&5;���bb�$Xpc��	^aWu���lgq��C�����&�"������{CS�-`��_I��b��e�@~�lԉ�7���w�ּ�>
-�4�FxuoP$�;?�0AE'˦��=�#�c�zJ/��O�BD;�W���2�e�)��$JCNa��[ّ��S�U�w��v�돺��l�%o%����O��\c$L�Q���AK��������m$ ��)�O��y�%��p�~7#*F���BT�]�D�[�����}/ru`۔M�����k���ß���b ����QO��jyF�&��S���_�un����a��NCwDT��?#s.�Ě�,H����6��&6S8��*1Z&�$�ʷ�{�H��V�jއǛ� $/�vj̶U�l���@4N%	U̟O���pkx��������3����h���g ʤ)�f4�����������8t��"[����GG���l���.ݽ��F'\?$w_.z(���v�@Ǆ%#�\f���N�lkrܷF�e�~~�MR�)��0?���5=�C#�jx/���mvz����m+�1��;qm�ؒ�a�E�ɽ1���?�n�t��rL���`�ԫ�M=hmFzId�/Ft[����H�:DFZw`���J3׊��/�o���"�=pbl�<�ݵ�!?�����]���3��"�+EN[uXS;Ǿh�=Z���ad�k�K<�>����q��G)�\��c��L�cw�7�Οw��^X�-2D��h6j�|Z`s�D�)1r��Jc��n�\�;EM�g���.��X�r������ϋ��������Gne[2�: �Շ.����B�@����ĉ#Kq���x4Vr������Q���N�v�"�v{� =�0�41^Z�m���o+́����~�����yZ���\�.�����6�ȥ�:���3Z�d�-[V)1|~���T|گ#��w������L��3&>�L[�fI��.��Z�(�H��(��T
����|��2XVb�q*�r�M��/E
i�a{ѷ����t��E��F$����vQ��5Եo��n��k��jA9�כk��W�j�8��>D�<�
��&�j"�"x�\�r,�1��,�����Zt^ݮj��C�����Tu	���!�@an]�2���?�l���3g& ��e:8A��u�*-g3��N��Y�b\_�+F���Z)ܸ{)�RrGw������)9�;� ��8�d������ð��T����T92�MPr�T��MA�������<b*����ˁ�у}��$$���+��DgM��KYix���&m���yЃ��Z�;���l3o+����Ӿ��-�A�|�2��@��-��5(a��;����x�E�D�G�:�<�X̱P�O{��;�%��9��o�_��X���� �3So���ClA4#ZȲp4%��	�(O�+z��@�����2!���8�����iL^U��FJ��
��'�O�����WG;�����06΍Mu[<�"�?
Q�E��]���`@LǪmJRY����){Ä��;�*F�/�*���LJ���z��k���Te	���b2�ñ.^�2R�ڔT�r�	a�9���_�Q3�ِ���Š�mk��8Z{%\9�G���&���}�%�}��n�a>�H��"-���cs�A��im{��W&��TjUT�����Q��_g`��/P}Ğw)VBuh������\8��'�ml�-�P��;��'fs4�c��3g�:N�]�Q>�|���]�yk�	>Jy=�e��p�Rh�v�1#^#��������\�'*�[W$V��x���Y�8��ը#���Db���1hg��8�	N��lQ$���f١�D=|���T�_ȅ��zՒ���tK'��C�oIIS�Ǽ������&�{�:W9�!m+��
'�kY^�7Խ�N_g�YnG��c��NfE�>��.��?�q��?��Q@�������D��I�g���нM1H�?p�����d�����F�{�vp��,n���6-d�K]�|��Q:�{���iѮ�ߒǢ�Mi��D�#'����e��>��2�㴈��!ZzU�g���2~(�{��,
 l�>I����p0*6T���>?��n-����zƻ�bZ�ӻ�ogZͧ�E?3bf��D[�|k�f�/-Wҩg�����r^�xi�_F�9��H��p4B;l ~������\�L�������5��B-R\����EƬX�N��)��O��o`4��ߠ<��yRA��E6�(/��W�Ի �q�sD�;g��6����1�16W�A�[����&�ׇ�)��w'���ݫv������2��ba�D�l��_'a3�L.)��ñO7%��|�s�d~�T�1�i!I�d��w_$��V�১�Y�e�-��:<&�aE-���U�Goʊ����=�XG����-�RoCE�+�/@��l� ��P��=��C�q�A����C�|ا���f���P,$3�����L�`V��NIt�p���ـO9r�j����4m�s���nY@$c!�S{d��xDlB�4�`�f�O�܏-�w�b,ͷ9������A:*�r�[:i�z�,�^L�+tz�X&�}g��߉D�޵�+�٢>�L�G���9�~��煇�L�LW^��/{!Ⱑt�_�*�Dƈ���.�a�d;65|�
��'��� ��{)��W�����W��tQ��C'R�f�d�i�
�*lQ^��a�ρ{����Z-&y8�����Y��F�={�${��B��5W�T60����l�O�n-3�!&2W�U���xQ�*Ӑ�1��b�����nө�V�>���^7FU�U�-�zL\�y�zư��D��Z�Cjp"�ԭ�VeY_�[.��r�	�P��H��A���|�b.8l�Z�g0Ʊo�L�wQ3��S���:�w  ��>jj2W�gߔU���̇�}��4����ɏ;�x@���]��r��.�=�]o0��
/ܕ�q��IG�S O���V2U���c^���\'�kx�U�2������CD^��������62x�(�xŞ~�#7i{ŋ���~��yD�V]È
��ԘN�����W'�Y�IkIL��o@g�,��5 h>OЊB=��6ܺ(���G�AP4ޣj|�O�o9�Ά�]H��\�ii�T ]A�g�s����I�%�����Y.j���� 2����C���W4K��m��rb!��ս�$6��Ձ(�D�
�hU�"l~�LaO��/����f��������v句@����9��d���k�W�� Y�EZ� O.�[�[tRu:�@�z6��+0JU��丗�QJ�� FQ�Y<�n�G��Is��sG6U� ����zȄ"�Ɖ�4޷�����W:X*K"v�~{u���H>�����K��V��Ը���*����Z/�K?N)a=��7w�0_�-(kKlж�L���~w4�ҡ�f<� 7J����@>0Z&p�gF>՞
Ri${}��S	%ML�[a�1��uB�����49���(��T��T�N����r�c�f�F@v�E�K���C�KH{x��^�	��]2+J�t���퐥"�+w$4rv��?�Д�>^Q�9�͝������:�����JGj��� >���sc��M�xgˮ����.Yf�u� 2u�'��}�Rh'���Q�a2�4v`�ˑ&�N�=FmD���~�2����f�+U�}��`ű��g7��P�]k����0p��V�0�`�מA5�^����M��d��(��(|�c�Y[*�z 8n���, A��/���;��:;*Y�Q�96��3�D-��4�?y�OGi�ĝs1֐=�00��7�}����qI�tOX�#grSƋ��F�D�G��p Lg�d���dS���T�z�R�[�+���T��d�s*,�(\�L���lR����W�-��ȍ��j�-�d@5���Vf�u�i�P����;�*۫���ފ #�E�R{�2i�Tt�^Ƿ���E�6� ��Q��:��σk�`�Gm���}Ҙ��4���	t;�JmR���٦-�,\����D-o��+����L%-6F�2�:f�i���+Zk@�X|��F �ӥ_V��>���]��	������7Uaq#����'zl�8NBR�:/'}�i�V��<B�]��es.2�G@%X�L��ҠI��~�z쑟�sR1��R�,ҏ����s�,����X�R�9L. -��m
=�O�D��>��$/E���W�Kq��,"Q2r-0 ��6Y�˽�������
���2�/+|�"���	8�Jmt|�K>��7�Օ�gA<T@zʆg[�~Q�hR��n>�=�d��muZQ5����s�}G�L] �U��>b��>����������&�^�҆�.�U��J94������
�p4>a�@p-U<L���CD}ظ]g��vQj��;��oO�F�pH��\����CuI	'��OXE��X���3��k+��*�Z���)*�Ҿ��T��#R(~�Fp�8e5	-�P���T���2:��/�@,���c&�
��W
.��Ӽ@&7���ZI��l�j߆jk�6;�9s��o��6 %��`c���Ћ�Ħ˕}�BU5�2�H��E:�K�A렰>4xm��4��_��|Q���`����%S���l�����u��*C��_oC{�ٌ����>F�V�y���=�$"b��	�����,�� ���up��C�n�/2Z������u9��8Ӟ�����:�BR��B-�D�h�I�( z���ܣK�+�0{J�5�ͤ�^S�����O'�}+,ע|����'��G@��5N�_��N�r���>���]��� ���E8�KBݺ��n��E�{�g�ZkBo�h|�FG�  �7������~�ա�G�T��K�������!�&p��;B5$L�)�Ax%�\I JA��G\�m�~���V��ZU�-ʺV�3����%9 g����Fއ1ym� @��\J�o�e�֝�� L�ؗB�析�Ǵ�li��cd�W�tuRD%��6<@14anN���F;۞��|���ǷON1 �W��D #HEmV�v�J.r���|��}���9y�'IhῇZa��`#���SM�c�,�7��)�Ə�gc8�o�`@��O���7,���=�]��mH�Gf�B��Ǜ>oX�Gq�06/��WE �A]ᅆ{�_cF��q��2�y�N*�k��x$�2�<���>���g�ѡ;<Ϻ��#���z�݂�rNѓ���_g.����q���w�{��'���u5���
zj��MY�����Ry2�+�L��^h���S@V�@�� v	���b%�� �QS��$�]:�o��!t�q�ͻk"�ԋ�+�̻7�0�h(�)7�Ȍ��O��dz�5��5�rFW~G���)+��?<r|3c��.B�T@�1i+�7D���BF'D 4Q;Q@�����l���w��x�C[/���3��vt�!1)�{��b�I=	#�yś	54Ȅn�:�-�.e�8�\��ʬ\�\t���<�6������
�To��8�z���ܻ^Z�a}7���
ŀc6'������%pXf!D?�c���ش�e����U��6
-���)r�����P��3%g��Έ�f�mv�d���.��Bf���ϊs�U�>��U:|o��YKl�J<Q���duK�ў%�`��D!�#�Y�e��UG��|+j
������H�0ߦ�UA��8G��'O�1��oz��}E�1uUp��5ɳ(���Gp-����0]�A���ͷq̼�]��0�һ���^��ZF���|�HG<���Á|���ǦY�p���d0�t�pV�|������"̏hd>�N�ˮF^�具�o,��O�(� fY���I̓��܇��)�3�^����}�[�>��g9���#�iH/��SF��������'���w��|z�Γ�J�Y�f��	������i����ج��(a.Yt�؅�	�a�	��4wkw-��5���ت����أL����a�	��/Hxn��M���4��Q����PU�����p�f�������㪶�,�XPLgv�k~�ZVw��� ��`����/���,��=B�kZ��gD��f)��zB��_����:��<Vr�gs�|j�^�i�sǧ>U�'I�ad�*=Ǣm���	}�8m��Y��o(������W����9�^ĕ~�<ܗ���̬�~<�% ��͋�����'Y���j�Bf�$�n!����o*Ƽl�gA����[�q�n���k����э�hjx�.���lfx��Џ��-`�/�҆���2EM�$s�3� B�|�^���韒"�N��3�U	r۞S�6T�IL@��h����R���ߔT"�V�ܟ���u�ŏk��MY��r�}]i
�uGVB���9�=�0MN�z��Z0��QT<APpF�*WR��L}��M�>OØ��+��F�D�
�\A%����I�d�#��:�.|��;�������̈́�A���~:S����h4F����m�f�9&Һ��z�<S_(�
u\�Q���dY
��� �
Sg��LV�q�<�������W�S�"U��_�M΢(���ƿ��S�]9�:ྺ�^NRF���c�'w��Ϭ��k�����Q"�2m[��7r��J�ھ������������hw��x�$��y��^���2� ���Z���$�7�h��Б�����P�=k3�O�9����F�W3{C�j���2pk��G�{?p}�S+P�:��	��p�"�n�g���w�!j��t(�5��w�M`�侀Lh�=b�� /b+Rϙ<�{�xe]���L��_q�nPI��Ϋ�v��D��G�Jq���7�P���� )���
���M�ҿQ��D��,��$���w���w�|�ڜ��c>����y���
Ҁp����΂O�[��C\�~� �f�1��F3�ǭEM�T���&[�L[����� P嗼��v������~��t ���[������Cݨ5z��Ve=ۣ栢�4Ѷ�(g���j+��Ma����[8�$��=�!�C����C���X�/z�/��+`���3>%�O�#���j�����)w;��8�H�7���ne�u^aNr1$'ӕ9�\5:�����{�P=�e\'�U�*�ğ��]���+]��p���ZFm�UW��l����5�"��ȹ}4�yZ%�H�'���p|\`����﷉�m�%��?}����s�_�xW�s\z
�dH��ܒ?a�(�2�;�n^��o]Kq��tb��$�����J�����5Y���=^�`G���r�ۥ�A����mӠ���d�����"�E�5|"�D'�������QmS���ȋ����/�3_����.s�ֹe����%�� R3?���6�;����ź��_���d�Ğa �{��3���K�}؊��'��|�y8�"o��ve�x�,�b|B~YVych��Gt=��Q�P�bBT7�}��n.יG����n)���PC�7�}6��~�DN����C|D(( @aq��si��b���� ����8X�U��U����50��Gz���6�,K+�V2?�8����\:�Z���5�L��8i��>r��X�32�������M�� ��/�z��5�w�C��C��Н�k��sX1���.;;����6B���91;>:�?-���M��8��#������d���Fu�I�H��R���[��h���>6#�O�����ذ�Z돃a�������R�d��p^��ߦ���R�`F���Gy2�RN7gd{�ʦ8X���;����ם�"�Wz�x(5��U\�����������hjw�|��
p����Z�l��x*��e���T�P����	��)��7$��V`�!�O0���\��3���ڽ׉/X����'@���}O�;�ҕQ�vV�\Sv���Yüʊ�8�S���[q�β��]$Q�]����6 4�ZJ�VHs�sa���M��c>E�˚��`�[%zCEY<�aA�W}$P!�����m�Ln����se�-ol�= Z���1l(4��.ـ"��q��!�$t��F]\%M�W(����~�k�A76��+�X�$�S�V���V�U�n�H��Q�]A����Ɔ�ۥ�K��S>H�,q��2���[%g�:�bء��oQğ*���i\%Ҡ��F���"ڍ{K�٪��|Y�z�Sv��U�+�p��mO ��v������ς�X���`"�-ҫ�8W���d��r^d�(h�"e�b�#Cbn�c�iU0�v}q����ek����pQ�C=�N; L4=�n�.-p=�"MS*ӽ V/���h�n���f��k�w��tˑ/��C6����+�sF�eի�44�fݢ���^�v�Q����MrF�%cZ'�-e��i�m��b^�\�w2k��dv6a����f��Z�R�I1���&�CB%��t.���M��I��Go+���W=�Uܞc=��o�Ns2YmS������ٿ�������ʽ3����s>�O���7��6�V�U�ܦZ&?����ђN�v�3n���ޜ'.H�C�- @gl�@�G1S��/cٯs�<
՗��"�a��2j{Ta+�S�}MU���K8�6�+�ph>�8oq`�5�9�q>n��T�nh.����['0�Q�o�[Q�"��� �o�dH��iBǪ�ޛ��7t|	�Y��*2������]|�}D_��)h���)r	t� ��n9|��^�kM����b[AHAS�<h?�$�e�����_^E���xRI�|�=:�K��'���ѭ���{'��7"�ys�A/��� <��:Ǵߣ�T���9����L���h�}$���ƴZn�J� ̂�������0E�d�3��ZojzW���;��L(y�h|�Д�8{�	^��Q<[s�@����k��P޶ہ� :�������k57$�6��j5�	q���M���R�ՙzr�`G�!�]ۛ��Cv/g�5U�f�z���dc���Q0������,q$�U��
w.���9t��ܹӡ��\�@S3�Mf[L��tªw0|���jZ�"�,�*�ʧ9��g���.ɷ'vE7�|x4'��=,C�Uqr3�=��J,��0���^�V�D��=nwQ�圵�P^�ӷѨ�^!A��X����j��'�0��)kP�8rhp��]I!Dl��z��ح>�����ֿ82��yi�~��g��{�R�Mu�p
�)vM��}���@�ޝ�ee���pc��l�Y���c�fbw!��]v9]�������vs�G�|�R�(�π��+���<	6xx

�̏���3IcE��U�s <��˞��" ,�v{�ROK���`M�9�/?}�,#3���5h���_��%�����DY~k:Қ���1���#V�wvF�(}-*0��b�f>�u��4d����0����.y s\D�FMK��-A1���q�V��^�H��S���q�(�-��xd��B�H�ظ���70��tkZP~j$�`�X��a_�~���y������J]����	���g��A�3y��g�t�A: �o޻��.E&��-�T5������<����&�~i7^������M��H��"�;���u�~����YA��M�ҝ��c$!&�j
U0��8�GF�=��d?"��S�91�^F�O7h�4��u�3�n��
"�7�>�'S�y�I�5,�օ*}�����S������7�s��]�2~���q�u�h�Iˇ��!�8^Ϩ���������v?�3�-�c)��g����v"�C�=��#"7
��cbf�6���:�mZM��ɷm�o����Ot%�m2��x z/�����_6��ŵ q�`F9 Q�i��}ÝpCO5�Н�w��@ ����ዬ���"&��+=��ʦU�K�$��V``�+�K���!+��4�j���2�<��\L�i���l���Y�c230`�ҝ)M�+AAǻ�OcB1��D��I��i$�����9�����B%���	4.>�(!o���J٩[;�p�qIzQ����Ν�}��&$4F�͋���pB��Dj��
'g�}�l�����l8#�#e=#�����(hs���執�Y��c��΁�e�0��J��q3��T�#�pfGQQ�'d�� ��;�B�T��+܈S�������h�f��/LO�nRq��K~�
`�����{Q�'}��W��A����n_A7�����+I�?�D�b82"�4Eqi�%_gI���q�"�����$�K�r�ؕ%9^�9�`�Z@sHk��D�g�FO�MІ�U��%�t�p}6�MLKy�"[�h�8�1���~�������9����� H�N�����B&����O+Z\r�J�W.^������Ge����R����;��Ԙx�v��ڪ�q���&��%�����>��i:��V�ݮ�d��]�������/%�g�L�`l�q�k3�F��z[����]��}�+\�Pj�Ĩ�Y�ȴ�f�`H�&_!۳�+w �T�Mp���%�)4٩W�2,g6a��mv.]O�� ���Hh��ɵ	��
9�e��(%���UvJ�|��������ju�6��Pؿ��]ϙ r��s��a�.�tS�#�L��J71C��jd�:Q"O-ظ� �29��m�/k�n��`#�RMNu����d�
L�x�iw���;dŜP^f��xθ��XI���֡Wx��zhB;/<"�6o�J;�O](��AO�j��~J]}��Q�'J�m��S�4�F��jņF�˱�L2c�|��t�AdB����58������'Ļ���4�A*�t�R�a
Eժ����a�S���-g	��Qk@;����7s�[�㈍k�."h�Q'�KOӂG����z��u�rQ�4�bbM�r�d�=��0Y�o����Ӧ�{���6L��_��٬�E��z�|����g�W��وg���n��7+��p�Z�����1�IZT�^�4rb.�a�M�@���0�j���W�$M{�Z���0kj-�1���fo$����NI�s���ac~�|�����gL7�)F y
#�N�r�,s
�h���4�}�v2��[V���F�4d��T�yİ4�i�Q�Γ�m@��u�h�>/!�W׍$v_�:�z�0��t�l��i;zn���1Q��m�q��]��r��]Ǉfi������|,��G���I�-������PrP��L�"��E]=��GЊ�v�˴}��ّ+�$ͲY�`�?�y���%���ـ5�2D� c
��S���j���h���G� 犼��|Ai� :ϳԘ6�����B��d��*be�+\�^�6�P����
Ȯ�DzwK"�}�߻+y;�Yh��P8�B��y������G�'�q�j��|V6�7��f=p* �>7Z5L��E�6�?>cIx�&��
x^C?���An@®�Ó�q�-?���f���"���<�LD�W��.^1XȈ\( ��v�3�����[E�#3'�֋s����k���մ捡t�%�����f�wnf|�pY?n�,#'>� ކ���)��M>��k�QYq2�N{��0د�����H�;� Wt� ��.�.��k�L�Xu=#s�
�Nr�5]#<��Jy����b�?�_�5Y6y7�H�Ea�ڦ�:���_+1�&�֕`����	�\�a4VE�ې�[�'��LM�Nm'1=9���kg�e�}Pi��u��N�a8���V��R�z�.4�9���piOy��,+�/1P�P��]-���/�Э8F��D�S��V�͗/�z��Ґb��'d ����t��v�7���x �)ªH�z�5F84��-�3��(�&�8e8 ��=��bU�w�D�����!�i����1�@y�W�&!Rx��2'�?$pS;�Ud���d��7������ˊ��f����Z1��������(�
�ԕ�r��O�x���>�K&��]��n�ͥ��W�"��м��==A�ٺ�)/9Z�n�޼3����K@����k�]�O��S�%߀��T�Zi�}�a��o%%����L��P�y�>껣��	}�v/ 9p^��/yςV_�̐0zIGu�j�]Dq�e�˔�S��N�8�6%�ЇHՏ��ˤ�D�d�P[�����-G��f�$�̈�k_؉���W�(!x]d	�W���V��5ُz�m�*U�UK��ɑ�����<e�'}S�p���Y|e-��bf��W�W]��e�S�ܸm���˖g��O�L�,c�+�_3n^�p����F����&5�Yd�!x� \���#�yQ�Ի�ʌc�C�I����L7�J�����+R?v��[��E����Ǵ����"�*�[�1�t����_�vó˲�$�v��Ōձ?�ޜv$���q��{��Ay�g�}��_J�T[��=�m�6���Z����ȍ������Yc�5|��B{h�76�#3�*�{��*��<�Fӹ%�qŊ�����$TYZB��$0��v���:�&S�+�C�~B�\T�^ϟ�������E��Ox�BVa�U�#y�/���B{�H&UkaҦ-z�z�]��C×Tu+����`��p�{��=D��/z���؞�C�It��M�Pj<���l��a�C�����U��G�'3Z�X�2S���'��,���(wD�Wv�u�9�bU-K�v/�葳�˶:�z{�����)t�9c���s�]oN|)�bH����������a�XÀ��t��b6��9��}� �^۰����yD��5��c��)<Ю��[���`ZJ'+���#�`�.P��\+q�����8O�傌�N����,h�u�p��t$��W'iv[�sb�~�)����b����etJ�0X�|���|S�,�5�ql��T%��C�]~��������2�»��3K��t�)��U�mU���:���jg�����{�z%�ۺ.~�2~��+�&�s8q��ۣ"K�[0L4m��Q��Qcg���W��V��2]��4� ��Svĩ="�-��7h�P���������^8gn҈
�B��݉yV�Y�N<�Gh][�����`��UiǀN�|�ݟ�=��´�������k}�9굖�.�-�ט�M;���AL{%e�8[����GE x�F�_��"b��`!���
���5�m�sp*_9^[)���&�hq��&�V �W�w�N�:΃�k�$��:��
�s�Ou�����>CMNf���m��LG�W���%s��i�c�W׷x���*+t�/�۫:D�lq6Ie�Jo{������Zۚ<�����<�Y��R��4=6,|�w l�w`snbD��ỏ�\�w��ڋj�x�C
)FM�u+��?��P�8h��7�%�K�K\	aMA��ĦҼ1�����A�� �A�C�]<4Ԑ�M��l������{�i����Y&b��LϒcI6t1�D��U�m(V�j��)�Ł��ѥ�w��
�E�r]�����M�w���	UyVU�����5�V��r��q����!�AF�4ᒴ N��*Ǌ�t�z���� �A-��z��0�P��:^(�?J?/gD�v���e�
'���P�d�oc����m'�(dE�ʸFg��z�(%i;QlʯHh>�s���	�Qs�k b
%�����u@^��F8�;z���M�G���D�OϷm!i	dH�;����%�1��i��!i��+K����h�{�*ۋ���d��A��Z34�~ƨ��7�����2ٶT�f�-�" a}�yg����`U�ⱕ��wn���kH��{i?a���iu��2]Plo�R�a��xTCU0P��������6��Q�eV6��+��z'���In��{U��k�k#�z U
�XΠjWT��(7\/|�vU�s׎�I��J�q��P�:�$�Ok�XE��1Gh�o6<xMJ（�e�b�aEΡ���U��FzW�e�"�!a�[�I�{�Rq�%�Y6��l͕=j֚W��CMU;���ڹ}2 &{]�r2�&�8�K*�4�1�w�������J|H�n����B�K�кB\���"(����{(k��kO�j�V3E���ܗ��u5��i5 A�i��� ��`�|�^��0��풝�տ{�}p���~�6���Et��(��p�o�������/��E@��V�那�x2�{&X~�
 �)=T�H�fU����dCPlT�0�cL�%��v��v��y��[���/P\+H��S`����+��/zԩ��ƚ<,�s�
�ލ�Eˀ魒9��	���F��D��a��&���s���Fx�����b�$�Qm �a���n���Y�G/���/�11IH�\�O�/�r+4�l�1��9�����T��Ij�Q��ECOcb
�K�#4������r0��:Ae���[2A��� CX���J�w�'�tğ���a��G�TG�ܒ΋��Yqz�T�:�~��az˔�F�[�KJ�Yc���ӭ%g6E܁r�{�����⸊�˗^� �Ʒ�xk���.Qf@��}2/ͪc8u������t���Y3@�tM'OX�te'9�*�a��%(H��k�S��G�,�̇��N����J� u9
 ��d��T�m:����T�KؘK�Ǎ	Q� �sm�)q�Ap�GB�m���l��iM�)��>7��F)
j�ߐ��`��%+�=�e�w��8p�U���3"�km#Xo���Ɂ9~$x��U����rc�JcJ�P&tz�J_lІ (�shZ��=��)��WJ����.|k������N��h�2�P҅3�
�D�U(�s�v�ur�uK�d�z��c�-�TI�����[�5�nVX��uj�����7���BO�]����� ?�S�"Fh1	ЪJ�Rd/'���Tc�Q	*�7�qM���[b9O�!࿲jr�aV���6�骮b*���(�f3VE!�Su���9�A���1-P���Bf��y~���]� �� �;�|��g��-�Q{�ؒ�n% �^l��hh�{z�)�S ���h7 fS�:!nx�އ�)��f/RMOǄ����;&N�1r�G�s7?��*A���`����W�&�� z�e��a�����`��^MJOnj��\��N��%�΂�a�������Α(|�r>��Y��vy�;��ɂ���͡ʫriqZ��q@ƛ+��@ j���}j���^`��NO��گ��/��j	��{��GW�/�\C7~���_�~�82�X���ko$��J$�w����, 9�.�;x��`;��6�Sy[CL�/wW&-�8���M��ݢu�
����6�>��"�n�n.St�kY�Ðs���'�kS�3nT��K��T�q��C���Yr�D��o�R�	�j~�9�C~A�\�'�VX;�#��?�-�O���@m������ǩ]O�E	�����Z��sY���{>��r�����7��Ϝe��� 0�B�S���Y�f�T���i�{�b���b~,n[����۸+�������p،Q�5�OX@K{��m�[9C�d���N�-ǅ�n�יXk"��,�iM�,�m�r�'L���Ln�`<\B���~|�*Unm�3^��� �a[�����N��ɲ�J���w^rբa�_�
f��f�����t _�3���j�؃d]�1eQ�b<��s��T������7���-��$��\pF��t�;�Ӏ�R�^��� �7���S�����b�M*��js��B�o�`��ۢ�2Ɯ[�G�	r����x4�A���TO-?��(�� ���T�CЭ�3p�����S���Z���kTkI�Յ)Dpg}�O�ҕ��s��\9�h���Q!��E�� _,Z׬�l,�y�!Zv9��H��C���o&V4�2���烅O��R�^u4�K�:	�(
���Էb�]r<v\�dc�V���E�m����;��mb��$���^ʃ>c�r��%sZ�V��[E#؜���X�\���Q�"��'p�/��HD�@m1=@2��.����S/%�Zҋ�m����4���>L_�u�)��|+�~ëBK�U
�;��c[���,�~�ۺ���}ݷ��K5UG��V�@A��O�}�f٦P�-�f��&�D:7�d��^v��
��ڱ7S�������l��X+�<�:B8�.�
��VT�����>�	sб3=�Y`����er2r�����٩�ߜHXٛ���aI�� ��rҳ'�#�mk��4����d[Y������s��IF��R&������|Boł��Տ�	>C�v&]+���"�v�SR��G�"ȝ��"�iF2���e'�͎�X¬�1~�9ד_
�@ؑ����h������Ψ����-^~+Qj�W��x-�5��d�D9㢁�����.ӟ��:ϵ�Y��b���'`��Rq�����m0���f}L�N7'
�
�Ȝ�� ���'-���JR"k��P<%ˆR��7�|('Zuo�fw���ޅ�Vo��$�qQ�nK�%
����x��c�e�]nά���SGv���>�DU��UU���+}?���m�Cb��U#�U4�Ej�� �7j� T&�4;n�%��ٲt�A���=���sR�ح����q;#v��'Y�"�n\엜.�Q7Q&R��X�-�L�3��֕}�a
��L�5K�W3/���<os�~T�KH׸�	Ye��!���y0}�P����Ɲ��O#N���d+fZ�B�4a*z�\�ʢԈ��i�Q���^M�]���S���� eS�FT PQ�t?,t��+���%:���sֻ`s�-��[�3�˄�Q�M��}ݟ�sf��ڧ9?p`A�h���Y�W�Y
�-����\����eq�]�׬d��5&<�O��k��!�df�c�Wf"�+t	���)lJ-�24�gt�B�x����l��­!j�-�o�߱M����C(���������� X�ъ>������%�Yĉ��L�x�j�I_�˚̇ H���'��
U��h��ww����~h7��-z4ͭ�M�Iz�䄤$i..�0mIu��`&NI��$�)2�A�
Y=��� �d��0e|�J�����ԉp��3 ���T���dm��ҀԲG�����o8`t�(Q�j������a�jDѐEve&g��
��#��_�5��}����t�.FJ�n� ��o�?���@ؾ ��;_�O�Z���.I͏�`�â3�V+�l�D�9���K�U3������f2M\sՓ���*�Y!˙F�j�T�� �t�����Z
A��KoK�!���8P�X�5 ��@"o��J���O�Z�v:+%��I����Go�j�*��;�+����s���8�?j��B:hX���+�6Ll\����c������$��(1�ēK_)Z�ǕvC�!~̨Qw�l�t\y����J`��-�Q��n�ܶ(��j��9�<K;�J=A�L����l�gXw���ri�'�kvBnBuS�
N�FYw=6�f�^Z�]H�-�<QPa����2���
�6�F<����D^iΐ�ȨX@Li9%9�?�D�ᑜm��{p��(��^.Î{��҂��<���kh��x�9#Z9��K5�a�����]�kE��8����a�9]4ڷ��_k����ƩXm��&/��n���"/[<�Jm�b��H-k~�n�Ok���{3 4��i@�8�Ԭg���$�(P�4�#a�E�
����������shu
J�A�դV_VOX������bx��趌�ʝ&DsOu�֕����0VJ0c�R���B�
��[�܎a�
�d��Pa喁VBkL��M�ٙ��0%�m�"��]���� �!L�}ƹsis�k�m���ҍ`Ŷ�����À��C���;����J�7��lO����ďՇ��`�k*ҷw�R�Jt;v�����&0���5���>@��Op.�Zqq��[�P���ʈ*�{�=�`�C�3�=��\]
1�N���]��!���n.�B�X�C��ьX�"���r�¶$�W��P����[�6�rR/����?���n�7��00}���Ȕpl/��;vZ��z4��٤�D�(�N�L]x��7@���ƛi���-)SZB��<N3	7��<�,<2<�N)�q�W=�r�"��I�0iP,��Њ���FyʹK�$�o:<Jȉ��PC��qY/���r�
#�|ЊB�]�6��*x���*!�y�6����'�kީ4��G���Y�g��Z*1���nvoC���Z���˫ �-ɍc�����xTG�hQ^��Z���q?� YL������C��N���C/a�)1�Z�(��������P�;����*�E"W�ރ�μI���E�G�gM nb����A�L�E%1� �I.*�(5f�B;R��GT[��zwԢ�����a����q��A�\2�)R�p:��Iy/�^Az��8��e�;|��2~��6~��=��k�P��A��Q��QQ�Wi��~��7����G�s���=�tԅf�{7���z{�]u�Md���xŽ�t\��k߮�2��2�U�����7#��l�(C� ���S�bE�8�� ���%��(ˍjp���῭Y������Zf� �m���@���l\���-"��ie��k��Ŀ��Q��SS�eX����U���6|E(���9��mE�\u]A�k (Y������EU����)��M���\m��3
q��[�G��+@#v�Ѷ~䢆,mu��o��y?%'��n�K�܈ډ5�oJV?���!r�8b�MT�%m"a�رZ����K��:"�.�a���rVE	+���䭳��"u�@gRM\��|�O��V�eaܪ�?����J�:	v�\=ޤ��ƨ�������(r<�J�΀��&hAЇ�e�z�hw���Y,CG!,�G˰P�����8f|^"={��� r�	Tj�� �{
�<n��ǁzD����R������Po������OĒ���ԩfGN�8)R���oS�1��0�z�u� m����^m���xRP9�;u辶��5\PZ���c��Z�9gEUg���PwZ]�>L���l��A^��]#�go�9yITI8h�0��d��r��` �̛����4��*|�5��)�^<u��b?��O)+���rF]L��� �&ݮP���~�>Y�v&#�l���y��i�IuN	��c^Es̬=M���~j�ԓ?�R´�.1oB$fg�9!�:U��~.���r�����!:3�<�9c>�\���p+F$����ǮO�o���ۤ�mKVuִ��eq��4T�X��w?��D�iKoU^���3�{D��wx������mp;@(��
�z�'j�����!>�@i��#?��Tn�bH�jRų�Fa�Y�� ��S��^H��p���b[Vs��ę�E���H~K�OA��:뮱�@z,���+��c�|���}R��?BX�����WRG8KԔ�<��$��S7�&���\�e���L����dxC�,o6q!���pa����1��la�����o��^�k�ү�9ÿu#!s4�C�����ɩ(yF��x2 �׏�
m�+�:K�uX=��`q�!�Ss�"Z���Tb���Cߨ��|Xt��ʻ`F8HK6��K�[�w��Nީ�8|E#�EK$���F<cwjDpM��D��G�|
���E����R�{A��:2��q(8��Z:�M��j��ɭ�ɦ������Я{{��;.�)R�RP��J
�Z��W�;l3ڙ��$�ϳH�B�\�75��D��+0��O�/�"�/��b8�F�3���#픳�K���l�j�ܦ���F�5� =�L'tc���k\� �W�_hA�
�0�4��pH]���d�{3�)_-�d_�b/��l��Z:5�U"y�d���&�(t����s���k�T�;Kw��k<=O��z�UG�#	#'q�a�F�+=SP��<f]tl�(ɺNqؗX��B������[a��[�Pf�ХJ>L!�o��� ���M(W��u��5��K�	�Q8X0qf�z�S��Ph7f����3��X���j����SX��f{򀡿�22�H�롼H8N�CW�Q����M�u��A7l�̑<�k�"�E#/ܳ��k��X��UJl�TW����4�G,����x��L��ؚƾ�o�
Pc��f�z:x��W�>̅���O���t��Ћ�W��i��UF���"K)����澾ޫ��!�3a���QW�`r���f�^�����r�5�=�B�(��h�RP���Q�Nx��w�c��B(s)��`�*���6�;	�r>!�1�� /u�tH���/;�i/���ƹ{���S#E;s��+厓�dd�v��u��hԿ�{Ɣ�l�(-�q[�� $k���U��f�^z�$
�r����Rh�)э.��QXN0̮���ț95j�\�ř�%��v�ӘFYғ,<��>_ɭi����6s2��N�ΕU��?n
ZB��\B߈ 1F�?�l��R(��K���˺�ƶ�'	nJ NB��M��p�a�J/�"�@g�p��x�7�I?�2�>:�)_���.�����8p�$�~ڸ����3Ġ��aBpQ�8���d��w��	8��,�p6�����@��aZ��](�x��`s���4Iq��JӘx��<[NT�b!��766ځm�6w��*7$����<n��Ɉ�z�u��ȶ��Cr�����^�;F�Đ�>�����++he�i'���_e�Z���[U��+ԋ�;cN���wڭ��# -�l8C�g��!s�+@��� �b�2|��l�y�A�Ѽ��"��u�,�|T������R��vl~n�����|�q��u�R�lа:���gn���&>"ZiL���v��	3�t�7�Y�v?BOmK�u*�Vg���Gʪ�H
4߼v��0z�&�����/��i��=t3�'|Wo�	tʒ
uq�$59m��w�4���!D;ӽ��D��?`��L�E��G���r�+M�O��E���.*���MݶЏ�����︤����Ko4�s�G�0l3��VG��MP�"-�L��k��Sb�7ɑ�T�)�&��l��}C�S��ʂA�I���)T�(t&�ZlF4��JV�Ȳ6���Sgkv�_B���kw?���r��ѱ�s棄a��h��5��n�K���d2+[��i� �<B�x�Y."{I�����pb8	Š�7κ��t4�!���C:��_�U���B=�ʌ���^υ�v����3�ci�o0���WB1+�:^8�O۴N�� ���G��%���(�F�?1'����ف���<�ȤIS��z�?��ݠ��sG�*v����~�����N�8{r�Y1N�w+�|�2a��n��L\�@�*Wؔ��n/�\S��A�׸���Gqס	��](([&Q�X�d9v�-�#�[�	�!̬Wߞ�fDU��=4n?���`�='����6:yt�}�z֮��5�Dep1�K��p�E��FU��oD�dj(J���Lβ��X�����h�>��<#��:��r��">�H=/�&8�L]�}ĺ���:�<�y�'	�[�Y�� �Ւ�3N���.>�.���e���'�@�U��Ξ��DіA�8KJ�&���8Ѱ $�^�9�m�`�s6�ܦ9�rK��
n�aHY�vJ��ޣ�FA��,����O����侶��{�bۧ�9%�@���,����D爵8�
T�{A���!n�R�/�'g�59y�p�;��y���QI�16mU��L�e�k�̦��m?�}��(j��ݖ}ˢ���',\j��=��lVV�[ܙ��+�,��A:m�>Y`�mUT��Ub H_�X�.[O��^b||�%Yg��	3Cxz�Jz�~37!����y8`X.��<][�*�����kV�G6	�!�8X�6=�[�:�)y���{����Yf���o��t�6s�ҵ�����BWm�tf3"� l7�T�}a�=� �D�N:Z�<m��Ǟ�`�Xra���E-rvhPm�˙��E�Ӄ���0KDY:�,��çY�)�P����L�E	�6� �+C1g?�诮,AyN��f&LB)�#|Rg���
�?;fًm�Gց5�B�b������:ɟ����rZ��[?�o>��*�Ǝ� ���0f���$�@0b��}9���b~Vё��c��W'��]T/���!z�}A{;w�.��
ςز�Ϯ�
_�9���:������S~�RԞ��3�S9Ǿ�wzM���_���������^I�'],�}�%����k����I`Hy�c�&7dDaU���m������O����1!�o@Y`�]���c�o����$l��Kx��+<�	+|��K�u�H�z�3�a�E)���t������ӵ�(hU����lnC�*v��A�
�۱��߃�0irbe�c�V�O���~T~b�v�|.�Wo�b�=�&a$S-��Tb2��K���E���v;�B�ڞMy�f�(�C%%l�����dۮX�C����2�=D|��M-���?.�Ab[��X���v���?,�8�|YIm�	�')��K"��`bT�=L��S�[��Z�ó��0'<3L����hm-R_�����j�))�r/^ <�<�̰���	z�l��ҁ�r&��F��B�P'6C{��XX��Q�pf�s��T="%�V���6�>9UW��+!�!t�/�R�ʍ2@�1&�m�9��.���g��L�vv�$ W'̻���y�

]�������߼L�}��`Kc�2Bk>(_Q�*3���V�_�ȏ�^XY�Ւ�]�������&�A�����ƑT�ni2jb�8/��$����̹�}�O�`55���a� �V:�_�2�0�H��f���"ߺը�?�r� ��.1����Y�U��Ia��M�G�@^���gT�rFW�3x`�C�k��-�TR֞�2�g!fn�R�Z���Y����y���Uig.d���w�-)��jw;��vO!q��L��ۙ�i
��k���E_?f���� V�7Q�0p|� �ܳG�I�v�(��r�u�l�Md,v�����ɴ;?��1OL
�A��= ��'���5��mF��i�7=�E](�N��!;�U@�&����O��%ݞ��q�O6U2G��4+�S���ҶX7�bI�ъ��HgrW�ݻ?8cG�ru2}�*u��
��P�)ق��~7a���vwi���`]o~uR����r��(����P� �s�N��x��u����[d?�'H�OW4��,���~�������ƒ�����oS��F4
{����F�����U�n����v��ԛJ:;}A=O�����?֑T���d��;�g�T���i�(l5��a��ô��4e��p|�*�hW�jOg��h�5�+��:TG�10���`�Z���j�5��)n��Y�w��@h!:*^j�{��E
��F�8�'���rU��-���ϻ��2�=�}7���A��cGsp5�}=Nר��:4 #�K&~Ք�d��5)�GBx����;�z׉9�Â	cN����)���- y���V�����zZk��*�<�`��r(g�(Ds���\;om.%g�GZ<�������HK��p�R�Ul��M�6s|��o�0�	�b��T�v�z��rs��s�M�ĵ�xB�"i�
c���aDF�Ɇ��'�e�Q�8[a�6�H�g���߆�@7߆���\.(�D���%��y�������%�Ze!�k��q�҂�	���T�%&8a]L����Oߥջ�FGz����h�S�DtK�!-xio�3����?b�N�+��l_U���TM%�36� �^���1up~T�	R������ŧA�}U��9��$�G���<C.~�/ġ�Ul�t��W�~5��D�|��K�RGkZS��x�Ӧ
J�"g$�ʸD�Z?��{��\���� ���`Rw[�4��oY�����D2̎���x�D����pm�6���,X�_��Ӡ�G�Rb�wvT�ܞ�Z,�ۙa����	4������ld�Pt����K'T��\�6OL`?˅4��}��ߜ�yǭt#+f$Sᬉ�Jz�Y�z���3|S:*�f�Q�p{���-��g�喳�zJ�OYk��(���2J�T��K��[��[j��͵���j�u�,kE��o�Ty���؄�s�>DnSn��8��N�w�|E�ՙ�um'����Q�'}�����4h�i��_U!�
�hkM˺���}��9��:cܔ���_{X7�W���Qw�3�\����C��A!m#�v�m�ƥ�$9D�"�{ �ˮ�t�q�<�w/���B,�)��<C;�H�nrݨ3��V�q��� ������)����B�Tض�X(��7�|�lTV{h["s/��DT�:2x%��>`/�'�-w��ޘ�J�U�����"�t^��#R����U���!U3R�g?��.utJ�۬%]VT��j ҹ����b_6~1a��U�}i�s���	_�!��^˪�B1Νɟ�oa�6�t!� 	M��Z`
ڕw�Y�Xk>z/�mAQkJ���%�:�eCGk�����<��m�ZlY�7�$'$#����B�s�	��YH��J
��<��R� ����H}PJٖ��2)��OY����"���f��=b�%������v���3����������b�0>�Ĳ�Zy�@�X����0D���^�n0���C��a����⃏Z�9s-�V&�����^A8 �_˃5cp8�q=뿶G��'I��C��Uy�1�ͨy�ԉ0`�̲ 	����,j2΄��_^�yh0��������3���?�)Q8� �B�wu�>tᢏ։�Kc���2N��,���6��Cȍ&7���◖f������	��͖u���#��N�5�pz�K|a�PI�t楎d���T�.�V �'(_��V��1%m�m.|�9^T�������xq)P؊W��n���-/�	ilm�9��y�y8�V� �F��p�r�ҵX�w�C ey����8���@���N��+�+e)w��?ȋmW����2Dp�{1����V�.d��i=K�^K̻��Ǳ��}l�0��UE�M*��y2�����n�O�9D�U=�4|oF]�[�)#]�~CRT?
m(��`No �tv*}2%o�,�@�s�.v?���Z���m�k�͑n~��X���U��Bن�"]�OR�F�Щ<�,Z��n��6���]55Sh���_uI�ϱ�3Y�d�&��MT�#c�zN�R(,���QW�c�����,����E�<upF��!c.������������a2������Ȃ-$��V�u���JU��!�I�������ܹ ��əc ӫsc���%� �>�I%m��1������� �mc�EV8��Xh`4�_�ɺ:,	�k�o'�l,��h�|�FM]��`��E����p�}�@�øU�1hDh�	�M��ϵG��W�֞��Ƹ�����<�XY�kᖬo����~�s�/?]��B�p��W����؁��h�&����v��������S4R|xhm�O�]4��ֶZ`��ń`s����C�-�~�iej/�2���NT�s�}���6��BIB�H-U�X_�E�B�����H�vּQ���*�s\ݣ� +���-�Yܲ�Q:��M�����z���P_������^�V{`�I�EG�^�]&Kh��~�9���t�-��c��.@�֐s��w��as\A9G!����+����DJ ��S�:�B��EZ��M�&�aѫҫ�|��Q'đQ����S{MM@5'B
�
�>��8, 3ЃW�t�����b,x�㤀m�Wc��xй"���%T�Tr��y1��RL9�nKB���U�b�g�_Zm(k�����8rԏ�q�}m��ͼ�0
H��G[M_����m]��{ؼ�1E�����g���W���.�1t<�}�DT�M�N=����<A��u��
�?���F§�	g�:�P�ȋܾ��*��u�nIм֑�Brz�M�e@��K�~854�,���1-I�}"xm�O��4��F�K��z��:k؂��M4���_F��MWʦ"��D�%P�����;���,�ֱ�Mv&�3?�(/�
\���j�o��y�j6I_�P\/����#Ɗ:�$�I���~}ߠ�o�l�?{@`eRc0)�
 4��S��b��I��Q��
�=z#�Y���B]�)�?07��*s��C��8 ���	9A�Ls�Hsh~�f5�G�j�^�2�h�f�Y��â�g�҃��0Y�U����ݟ�6�
���h���~^��[�@q��ֺ�OU�~5��_���=�E7!?���x݅�@�	_3� �~Y����nة?�Z����YaJ�MIN�$rv���v��[C�ڤ��)�����B�m��J(&!��^�+��OHg�#�h�6��Cc\�r��d�=oj��P��vD�\8]?�wAr�U �j��| �/B�8}-���t����t�4�{�!g0�����C��%+F�E�D�+�'�h�P�(2���AC+���@��/E��������G:o~���a����
�|z� �N\t,� ׈��/��qC��ђYoф�g�J�DF9�A���"|��jg�� �w�zS�~y0���ZAja2D·O��׊J�z\��'w��$�Lv�7��ۜv�^ڴyҧ�S^��G8��SI{�Pb�v+�[d�|��ʒf�ٰ�^�ȭ�Jo�� �U)pk�Q�����6z�aU��f��n�z􅃮�6�Պ�Oh+�-|*�<��G��r��X"r�V,W�ە-C;ǗC֍��?b``�H\5F��3�h�`S5���4:�@Q�-�������h�{*Y�����k��b�7���O��߼m���y�F.d(�2q���q��� �9�h�3�Kb�߰���:ZUr�s�FW�c�/�F �m�� �CQ��G>O��u<�B�ږDw6~���cp�SHk3�X�X+�<}x9?~ �*�%��#�+�g?
ShS	�	�#��	���B�V�0;���8���U��W����O��L8��h�y
}܇�$	|�`tX_>^�������skZ���t�k��kR������R-��������ܪ���F����gfX;�~U����Z	�s�J���%8�SpS3��7/���W_��vA��n����Y3��65��B�;��v�൲�Hw6qvpJ��Fe$�gQ��A�������R5�ҜJ��}W����d=�莪��!t�'����� �`�k=�i�r�?��0��u
�ZL {±|��(�O�,�L��y��*��P�8��գ�!f��32�Z���Yj�y��*���+?t�o�7{�y��������<?_�5\3���{ۇ�#p��si�8_8r���M���`� !T����I�dgɂΔ$F� i_�� IM�&�L�\Gq�P8|ֱʙsM�J]��R]u�i���R$kj�Յ[�w�/Aɩ��@sCrC`U����<�UHzj9����&�ٷ�>GY)��wc ���ŭ����V��r�Ч+oC��Ī�K�u5ˏ��I�T�a>���f4�s����1mG�0���4���C�s��c��m}�X��|�
�99L�3�r�"�$��YӐ6�#��g�aQ&���r�`遰�]d�P�t���aA�F(�r��Jb0U=��ɜ���X}��|�H&�i�����X8�~\�um\�./&`��訬PX
�zb���^c����ϟ�ˊ؊8U3"�-�G�r�v�\"}o�����<*h���;zGR��`J�.�V���ϥ��dH���؄U������۳��+Y
o����x����Z+
�:��wg�Q��i�����)fOd_C�e��c	��?��%�r�j�i�J�u���8��B˙	�LY8òyڳ1m{��V�yQ�Spz"���P�^H�ȝ��x�Ii�>	A}��
"YR%|�D+{!���ap�l����^͘��h��r����bp�jNG�������s����d�n��R�{�Q&5�dbb���D:����WZK g�{j�L����!e}<��7�q��v��mԸ+�?��gf<��Y�`����9�\�	�eT�)63�j*�b��\M=N�:�	���֚{�;�p��J��\���s\�X��`�q�v���z���|l��yLXK�n��P�DT���7�����#"��N�
`���^V�E�S�˥@`�{��M�+��L�>7y�cAY�&!c�V��I����F���~{���G���;�������:7��V������$w������;0Vn�P���JS�(�H��Ⱥz՞�w�'�`��W���Է���9�6��1(%S�q](1,��A�����E�I����:o*&JR���h����r�)1ȟ��\��?��=Ԯ�O���!��
6D���ѯT���sU�r>)n��US{�e1���j_�)�t�El��Z�?�oGiy�\���W�;�V�/�0���6l���˥�w�l��R1'����,�r�.&�F��������Ön�
��#��/9H�e�X�Bb!
�qg���m�6��K�]ߓѐ�r��F:gI�m���w;	��u	jl����4�L	���q�환W0�n��_a�]= ��;�{cRЂ|�/��,�֤��+�i��|w����_��m�H^�G��"�"�i�Ns�D.C7�W�=:�O&�<�����4e��3��t?l���e�L7�_=�*/T�����<.9{��oG����8KX���$�a�k����<w�Y����՜��k�G��U�X��]k�il���X�z~����:�n�U��Ǩ"����8���ì9����J����q.=���ѫ�9I��=�5�۾�$Eu�w8���F���>o=	�ε�FzD:�[��,�O{ו�(�j�S~C4��@��`�m&��8k��V����%p�ά��Sn&U6�����X�*n|�B�tmʋO���U^�?�8Z0Iv��P��g�$Ƕo�qӂ��{c5^�Z����3kf�YU��5��ˁ�[ K����O"-��zwW���d:$�i�^F�Xt?�,~�lYM�~�?��� Y�LR��}Ψ�0	"���m���9 J|Ll�f�F��
Ts��'.n=ˠ>�����*4̂��x�c{��2H�	f�L�<���rU��]x-,+M�ig�p|�EK���Ĝa8��fI����5���}>d�k��(dG�$���y��tZ���z�����ORH6Q�> {҃�H#я&@��(ÿ�۴B] ]rƬ���%*��z��@o�t����D�Zh_�,���<A�ӵ�Y�����\���ث`�����t]������3��~���8�#yW��a��wUVÓ�4)nQLrˊԡ��E���MM��7f�����j�BێWc�#�G\�.�C6p �1��ݿT\��`P�n��7ܔ�"`ڇ�,��ײ�!u*N-:��~�"�K-���7�&�`���5tm7dQofJ�`�3��Q��w6��
�ڿ�X���v4�RJ4v�ߺZ�#r#reg`6��o|���)�����O	7ozS�7�*Ԍ`Xw2}�o�d�j6�hn�[�����Z]ɋ�Bv�^�G�EX�S1�M���N��G�e)v��xuM�K������A���_��+�� (l����g��'���@5��ݕss`��Q,���D?_�!(F�E`M��^#qS����`}�Z�[�"|�(:@��1����Ӓ����,ɹ��[X�-�
&F�0��ە5ܢU�wa�)ô�c��:�_]wy�����p&��r@���'i!���8�%S�41'x9��D���^�䴼��D�c�����ߔ�C���nU��)n�NvL�(p��b��������-�l|
/ğ<�����'��XMP-(k���ݱ�<�3�m2�4q���kթt�+��a�>P�qUlH�y���\��p���?ݳ�C�9�7�[`U��M�z�+�s�wU��Z8/8Qd��Bذ�\�\�0ʅ�NH�b<���*ts����C���y����{Ug��f'�)��黬u��Xs7�#��
��8���S�%���R�����^�F4e�ߥ������0�h��|�_]��7h��'�ځ��f2�9�Z����H<,Z��^�S��F�u��>�rr���u�y+y�r�����-+Ƶ�
��^�t����u��N�~�`�Ǚ80<��Q���Ĩ�+��ZJ��_���0����w��	Ei)j*s""_w��{#����/����H]PIqˢ�r�_S���"�޶�;�6Q����g��Ĥ+uꉧS�n����d.��h\�Q��#
��ܘ۩<*2�p(D+�B�-W9U*�p�Va����^���ʤ��|e�{���yͥ3kl#1Zq�Bn1�)���$ŤK��9X��T���p�{5�k�(êi�PG�Q�J~}.�^L�b�pI�T��lMﹼbd���f7�����D�L�qF+9'2S
��i?c�k;�B	0Ͱ�5���(����gd��?M۱��
���*�_ʂ���!��D��&�+�s+�����
 ���ud����'خ�c�*�K|��bmomYr���H�i�T(V��4߄�z�U4�b�x�^�m�㇍�~E=1Qf�C���%��(&q�|y�4t�#�k�XM��;68�Q%��9��t���~J���l&�>��k�[sun/2��k��c{�s��߬�h���Pˑ\ u{��U��ٟ!�~��@��8mA\�s�/�{��:�s�?D�BNO�E8�	�Z�*\
�|C�w�IF�G��b�!�`���1m��FXnR,M�3"���t&㋚)���Rd}�����j�b9� ۳��#�����I�ҎC��ܘ������m�%���?Ϯ�V4��!閃��@F����:BM��\����p�����'_���TH���%?Eë< YlKM�ՇTD%��	y�\�>�:�t�:e�o�~��V�#i�{��va����2�f��T�(��%��hh�s[� �cy~@j�H�7Ά��/�e�=��(f���R�@^#V/����i"#aᯕ�Wp���ѯ����J�MܕxˉF������g+�� ��9%������e��b��u7��^\�%A7�q^��'P�7���wYl�������w�h�v�ߪD��oC�4[�!��ڮ��I�35�C�C����ϴ�y���R���'[�#"96{�_����U��x�>JϘ��YQ�;�.Ca%��-��t�d��Ɣ�T�B�蟏Y���ΈX�auz�q����b��A�d���x嫜�u	U��+$� ݝ��z�n�<�]��wS����J��#L�5���0�Y��t�G��)|�5�]�x{}ǋ_�^Q�l�w���47��q9�h��A��	�>:J}�/�����Ct�K�IV�<̪@��.H���q۔I�nX�W��0h���BO��k���B�@r��y�*ZlDN��(�/�G�I`��5׿ؙ�>�?�'@=.}YsT��e?4�
���,Hh�gs
>����^Z��xUX��)f�2e�*Q���� ?V%�e��=`� ���@Q����f"�K(K6��8�LV�vPG��qS��2�n,�u���4k.���c���#ʽ�(�:ə�VH��;<�N�]�
;CR�A?;V��.����1N�qc�!�m?Q�R� ��	h6b�Cڴ|6E�W9�y��	����FCy�az�Ѹ�q������Ժ��!Ea���;'IQ��;?�x#3����E��)=rw�֤��O����4q� �o`�4��穨u{�_ȓp�ݬe?��B��j�E9�'*J��pN�:�^�)��AzB'�)f�8%�;0���)��f�	e�YK�>6�侔CF3�0�=>t
� f$�B�1�$Ț�Y
Hv��(�z�o��a�_��I��|����IB�M�$���9��[�*Z9�ð���晸/�Y؞7�<��:Z�F0��I�>�IJ�����݀a��8��7��*���
Ԫ��t��[�$g4��~w�%�P�JX�m�3���i~�ap��Ϛ�Uk����o�|���k�0�w�p�J��C��P�|<,�uIY���홻a9h�i����2���Y���^�x�`�j:���T�4���%�k�ڂU]��ᛖXW?��DƅEi���;��Q+�:��n���`��r)��g0��yƨ��?+��n����-F�G}����}OU����g�5�Ma�'(~�ґ��JC�	�H�+����k��U�b��<?	�`s-Ǫ}"�ӧ0���C.UE{��+��J����������t���!�L�����X7��&m��z�O�,�~�g����)\���X�Tr�̖W��=��Bu�n��[ �U�=Sc'.2�f�U��m2�W�nߓ=u��&��E�4wg�i��%K_ov�b�o(�=��k�� Җ®��	o��X����	����Eu��;���'w�go�B*�H��AFxA�FW/�yN���@mG!�\W����]_'O��nٷ�@�G2@�����a�&�|4�1�����������<h�D$(�V�h���SK͑�9�W��C��z,��2:��2�/$)k���Y�G�"S��/ܿ�h�2�u�iq�6�>n���H�Jv��>/2)��hp|rǺY�B!T��L����u��{��X5o[�h�|�� ��N����x���2���Az>po�3�eP�E����I]��SW�ۅBAD6#̉��_�l9Z��6N?翟�W��Ь�lQ�[�|kD1��cd��ɡ��,)�F��z'>�YqO�L������^�t�:`��s'E�i��r��
�xX��AL$f��<#�n����}-pf`-7c$��h~�2ǣ�^i4c�F{{��Ax�4�[E��(Z��ocn0fQ7�d*=˨�!�U姯��c�2;�C�ѓ�j�(�b�V����^�[�$���:��j�:k6t9���e.��.͘3�h��!ٽR�5��OZ��opr�>f·S�O{�Bn��ޗ�����k y�sB{�,p�_�`v�s)���2��b]�����)�+��n�1�K�����!>�Ԛc��'ol��\�t/V�g%���i�7��)��T��V�܁�rRH�3����ά�����x�ʑ�Be�%�|'�#��T����jR�i��$IP:����-��cXS�+����	��t�\�IX��|'J1)�`����ar�F�f�R�_姏������u������&A�J��?q�v�?�}�Hn+_�d�:{#��P[��cy�qm��h�"&�]��s��jX�	I1��+ݶ��\i5��j(o��<��A�_,]v�J(e�& ��b����%vb�ɪ���$U�IZ3y��h���,���v��HLm�BrjW"�v\t,�R&1�5�.h��ތ��-o�_�X�
FV���y�^k�X�X��xB�u�[ +�V/Gŉ�ÿ��[/��HWC�&KΑ�=�������
��,���j��̚eMfRם?LJ���MkŦ�ڡ�+ǝ`�8�3�Gr�Z�I�V� o�i�b�����'��7�+F�\�L*ϖB���B]B��yH�$�]e�y��S	 �B��疑/�kI���<�E�hw��p��w���C�w����C:<EIL���d;s%�b��;�t��Hq&�0�;@��6���M�*3��&�A9I�}��ܞ�\6�UN*w��?Vkfᜥ�J���9㑁^��C@f_VU�3�n�ne�(+����$A��-	X��]�I#��e}�1Jm��G�fܚXb�y��H���waL��]ZΕ�,��:5���^�dl阝akM�ǐ��Yu{�ļ��J$Ce����U���]f�&$δ�V��$}'H�X�p��Y���� �iͼ�H�J1R�3aZ�l�Z��c/�w���D�)I�Z�����j�LqN$�W�[�>�V��	g��u�2�u-O�GF�@�������kP��dZ>Z��`�w�*�6U�K��"�k��:��K}��QT��˒*5�#�(���6��<�Q�X��`�!�۷�)%�l!y�<��I�d[b��i8�~���JYYx�Q�a���q����Hh	��jF 춨7�Tiеm�)�8��]he���F�X�n�y��U����;�މ��6d1I��4 �E������2Q^��cI��Қ���혇5c�Ɓ	v\^!c�GtV�����wz��� F�/�c�����%BV^��̿��g!�^�(��v�����qV��1�Ǧ�QƂ��,�q%g�|�m^��!>(�gd!��x���>�F/V}yi7K��Xn<�Y7}>}� �����d�m5��
wD����t7v"���h|�C�{�kOd7��ǛO�+�?�"�6%*�c�R8C4�*mP�}��סƒR�ݓ��x�M$�S -���љ�T�F�{rզ�k�$��'Z����j������Dr�ɇ�v��
'�-I�E��es�"+���8����ܞ�Gz#7�����x����=��4u���O�'��o/���20#�c�:�qgxy�NqX.u���"��Y��PIk!�-���T��?�+�Y�M�~
�	H��<f�~6P�/�M��%c�ՏD�aՎ_G�p���xĮ|�46Mg�v9�;��eI�|�Pvco$0>��i�Q�
|.�jˇZG��E���a���˲\u>b�-㍌��9�F�,��uԷgSB��]�;��#Ё0�JX��q4[׷�܆�:���sq�6��1��<�^K�&K*}������v�-aX��d/� �}w����ڝ?��cXwaOn��W�X��F�����k�ep��ly����Ŀ� v�yb�yP����5\�X=R���`�E2��h
l���mgc�b�`]�\�J�!~��n��k��Պ���Hjs3�I���d�B�+��U�����W�̈́1ۆ���<2��w�[wCTVn��(�"A��u�GR��*�j�}��1n�e.�[a�����'�[(�Ø��hi���K8��|�K����v��ώz6�[ʍ?��o2��F�E�*���-�vgQ����&��HX9�1��5Џ���8<�BH��vuG���&�3C�j���H܄���봹W7*��%1��9�����2YS(�녨k���oᛛk�f���A[7$(�\�^�z��r/�&�?�F�����je��-P`^��Xq:ɥ�ۺi�s��C�п��}���Ň�O��,]����=d�O)�q�S,�yf���5?G���L�?{�*iS1���Mq�2���:����Ă�c�pz��	Z� ��fR�%��Ԃ��~�����	zd��($�w�t�@��b@+�뎲V�wN�6*��1�U;$�����ٕ�]��ia�⸙ gۊ=>�S�ÜTmؼ��dȽ��?���u��1����_	�g҆^$��+�����}��:H�!�)��1��+�0�m@M��T+�i��i�aY��nf���(���j�6��3��x��!�g0EvT��l�V��)��Ԉ b�ը),��t�ǎЦ"8T��]]�i��h�l���,<Sj�z��+�ғvƘ7X$�����ef��P�uul\�(�@��bv����yq�z�����10��;Gz��E
8�-d�I�e�e�WHL8&}|����7���5�9�:��NB�N%������� \u�|�02.#9#t�������%��YS�e���>�P,�E�ʾЬ���c�Q#Ȱ����xa<�'0�+�����T�[��c����^���'��^.V��#�A.o����T#-�9�~�Y Zw���}�G�G�Fcx.P�m��Lʹ3H��#zA�Зr?�A�%d50�D�Iz/��}�vFj����t:���QL�����bۚ��׹ݮ��b]Q$���2�ٽ�o�����g�+��5���7�.��ڻ��J{�q'���^��@��e�0����7���r5G�gm�Ǉ����[(ݴj~���/B���R�/▔9�������
<�0?�d$��xA`@.7�8���V��!��SW5�VW�:kd�:\��Wf	I��Xqss��h��p�@@`�j�`���v_7��
᳑�������������[W�zz�nu��㡮�������;B��v�j�r����>���3U,�����?=[G��	�-�Okar��@Ɯ���]̗RJ���)���f��$��1��PB8�i�:!g��Q�a�[II{!�j��p��%'�~.��p�t�o�rT��_�{փ�&�%�-!�i�_�
㐇���{f��!�8cT:���������z��KӦ�����J4��ܸb�/ڊ�h�h�e��Ub6)�SE�f��k�bw�w}�M��2Cv�"A&"��M3_/��Û�����`��o�}���U����ެ�~�?��ҋ�ˎ��H���+�!6�cZ�]�A�G���oy���Q��)��Q4�h~e5�xp���A�o34�1v$T��˲^ w��=����Â���D/�@�p��>�b�f�A��	wVaU�ı��T�ƴ� )`,'_�v)g�'�
1�ĺ^p�~,�x]?����a7[�'ur�j�Z�L+_�xo�$�%���* ]g������t�Ϭ�/ֽ�B �#�!H�|�����	��'s���rvwG�F�۸L�g���h��.�q�3W�=�#�� EO�1��;{*����<����I６�y�oж�E���~T�\+*͵B36�����7؜o�S��PŌ���%��c��n��I�n�k214ԃo�N����0��(=JE�ȗ���y`O�W��g� �6��Ź��ٷ�x�[���k��Uc�­�ejqQ���|-�ʊ)F��l0s��(�6�
���!�K6�`��c�����rb�R���ܪ!�C8Mƪg,vK�m`�9�>�r�J�)T�ǣx�,�HtZ#�&9,���P�����yf�����^�����Wf��� � N��*�܇N����bҒq�s�
��v�gשڲw�q�^v��Z��zb#'n��ke&��GN��4��I�7a�)$4�@�<t�̂�0�o����1��^\���g���DH'� E!4��Js��`�A8��r���;��GAG�V��#"-鴨�}3}V��z��N����M�ݪ
��=�֑�m
��o�fNQ��P�����L���p�bn�y",ř!U���'�9�}��B�d�@a|2Ku9մc t�"��=�b9��M���öX�&Vyް���X[QE�!jb�ȷ�"[u8����_l�/���T�p�OXԸU;Q���e�wu�������.�l���`��9T�r�Ч��q�C�!�]�-�=��4�_���q�k%���Y׃5x)�H�.�������{��y�|H&����b8ͷߋ�v[Ճ�)�$Q^ڧ]�Jb����W&-�`\�|s*���
y�k��%�ܡO�7>�:덞h
1�P��������I4������gK �Y+p ��k������V��ňt��\�%����\֞�wz0�B�g�EZFq#c�xZk �j���H ԅ'��}I$�R�h���U5�/��8����1�:�0IO�OU4M�Wڐ^T	�l������No�e0�& ��3�ǬC��.N^�$7Ck��3�!4<a@ ���gj����6p���l)qlb�+�C����k���R��%mDBiM�3�����80��Jv�(��>W{�Op;�aJ
E����q��:����?bgLp�Y��/��k�8EV/�m�"���w�Җ��\�1�<"V�ɺ(
A��V	n��\ �m6*J�1����E#�#=�'�W�(���`�������S	
��$��X���"������;r�%F�g�M�pN��G,g�{�H�PZ�\9t
꽫���ܚ�|Xv��u_���݆�l:'�q���)���\�K�:t|���~ �uN��SQ�=�3Zr��V+�塧��i���;0��X�nTҧ��{@�͞@�����L��v��ˁ�U����K��=Z׊�y.�D�4�OJ��C{�^D2���{݁�׊��| ��V�Rh�--�����%�+��C���Z��aV7�U9k_h�2+1q�#���H�s��d,�I��6 �b>x�����a��nh����u����j�U⼹�v���h�V�ƕ�JE9��G�j�	���exb�i�I��F��t���W�g���R�N��U �%��ВƬ��Pˇy�%���dY�-��@�(��j�'������!�V�i�Y[bT��#�B8�N����7$jք*=VR`1ITa�2=��l|l?N�ωIFFȴu������ZBg�@�x��`&)���9\\����!!i%m/*��ߍ�*m_!y�T6P<o�H�FR�w�3���5E�g$t@���\m�F('f�����!��`�5��#��aj���mH�R͎�FT �+�aY���GS|�nݗ�⿆�ΔHc���4UGN�CIN�+/Cj1T3jU#I�ς\��<�
�(�*%ln�`�ffX��<��g�AՐ�T��)�E>�]f�N�4�L��t����˔i�~B$�~�hS�&����]7��eKx�E�i�݂g!�I~�[�e3Qs�F�����	�Yxܔ7UM�'�v���!uF� �+��I$�j&>�G���)\.��*]'�?�R�"v�$�X��͘�V�;�A����+��p��	XJ����@�^���ʋĽ��eW�w�ߔ��v��*���*塛���IzUGǂ$|E�9lݥ���+
u��s����gXj�_Qi�j�z��)��sZ��]0�#����ˈc���qM�2�І��_;]Yg�ߓI%�S���j�D�iK����?��aI/���
��	?
��t؃��
��6�~�p���3pA�a�-�~��^��@�
Q`WN�Av��?��R'�D����XM�[��٧
�r%��OC�Ђ�1��>�yfpRw>E��P��P�_I��zB 7��z7�Np�X^�ߙ�*�d�]�o��}C��WDbB�ϸ!y�#�E*bž��=��eF�8����s�w�Uf�/�bR����B~�ݱ�}�s�S	܂E���P��\�����Z����/�/�?F���Y�1����s����uևI���X=��[�x A|��~�4�R��oڧf��o���1��I R`�������0O��{��-d�o�4p�7}��x�˸�( �+7����g��Ȍ�j#B�2B�} E;�T�Кv'�ژyn��Q����}l��?���|�׬\:`@-���l�	�g7�h2Fjh\vX��v��z�$��:�B�\�ۄP��HPB�������fC)��7�+���a��\����>h����PJ����{o[3C��B�?miWwV#����z {O�{�	���[���u����(���9$P�g��(�[L"]P$���o�5��j�ie!��!촔�B�ĥ���;Bm##����+ɹ�Vae�e� 
ｳ!/PF)�8-s����2�7���W6�8���ԇ�zn��p���	X�Y�}�IQ��z�#��Y����2$�X?�>ּ��Y�E�ڍ�{`�z��S�ڋ-K��5#�H8�c�@�8ʌ�jg��]��"1���5������o$9�%�*G���<9�ɏ����:Wwat�jj��'��`H�j��Psh{et���G1�'B�����a��7O�A���G��K��2�Є��BZ�±�Ҍ������/*4�B����	����Tf����3�;Q��	�o�j@��&�(~�T}�@�5��qj�5���1:!�܈�L!g��7N���I���KXF4��_Âz-f�����T ��VwԳ;埗��e�gRDM��!�w��+%>O��o^��!3�b�9�~�bs�7��s��*�hV�~ص�i�������|{�C��.1 {��5Y!��}�b����랿�s�͑�No�Ą?bs�H۲u1]�ըc	���I�)�:��	�N~����q�ꅏ��f�lhi+��ғSvU=�0C߷{��-s�r��Aq��}<�Eh}�/�}٤{���+��ɐ�*}��h ��5yQ�����Ƽ.@��9�B2
~��D�}/N�t�V`X�R�֯k$SW)��eZ��(ҟ
���%�A���gx���|j��
���u�b-���Ok*f����%J�wu}O�}��&ܧkc�:�P0]�"8}v��F]b���e옄<�&6�M�k��,��]��g�� c��SF7����x/����)�I���X#s����,���Ô%�UIݍ�^��n,�7S��v�j5��U��x�Y^T�Zv|'V��đu��"�(��}�Z´�����ב
�5����D��*A�y��đ)k
[%pn�����f��u���=�g�fEH�������*�O��q�=jJ=��Gܝ,?��<
T`[�������w�YT��7��H���Δ�I�e��I�G<�m��I�����Dƨ ���l(���50��rmz�w^e�z�ި+=聗_�� ���}�Zf6�fW�F::�>@s&,����R�pOOu��}�Tx��BI����G5�%�4�+>Ñg�/f9yJ�d}��C����x�M��/X�ڷQ?ut�}�O����Ҫ9{?��㻿WA���tMl gdҸ#	9�=�z�;�jjb@g8�@0��#?��4�̬ab?�45�H���SkS('�Xq�}�;�@�Нk��y R~���$bu��p#C�R�]�������F��@�������ՐN�cz�� {�4�+	��8#��S����s��1��SH�i��
��2T�q�p�|$�w���5!o�g�K/o"y�D���<����T/"GtHtV]��ޡh�|
t޶��Z�Ww���F��[s�qBԦ�C�	��~Ros a�
�Q�\�B���gc��io%2r�^ �ɻ#�^������1��lϺ�حs44�/�	��9R���N�2��!�����Ё�`�<���dӞ���I�Y�n��AQL .M�/t�pZ�*�Dƺ��sq�ԧ��̉|Y��\pX�{�j��R����@����ޡ�fs5e�M�\�:΂��C<\E�Z�B�,�"�B��KB�5)����F�[R���9R��P�I�i�D}�����n����Unr�PʺZq��39oY�!#����o<��E�4p#D���:b���F�Ԇ9v�u:b�Y1��$�U�	�&e����_�
�fo��{+?�S)Kst+Э�.�]E"��r�F�'�5���F�H�'Ė��o�	)�`�d�N��Y�|�q<P�o o�z�A+S��q�I4{�&Q�	7����0�j��2x�c���[�t,���[�q�
"�KLڏ5�ɏ��PǇ���f�=�R�
(��I�8¸�*��n(G�''Vk��M5�rd#��[���";X!3Q*?!`5DЙ�+�� �Sz�8��*B�3q��˓�=H	��^B�����S�x+���|{o{�#[j:Ϯ�p�i�}�^ɼ^��OR�#Ry���p�@�8!X��m�-�y�3Y�(Ʊu���`�m�u%�p��+�&L�&r@����7��i]�T���7���=��Zz�y (>����%0(䅂�5��N��t�l�ȁя8�i��(.5�u� Ƚ��O
���%I;�x���dx
�k 2jY��
��΃&a�\����%)��x>+H���/P%M:�x���+��U!�i0�z�p��T�o�����q4r!ǳ�JNsu�#�CYه'�r�xp��uҺo�����%���A���5Y���CS MWkª函n�f3È8�XyV�%��Y0�%є�h���4�	f/䢠d���h�(��?����qe��esm�S�M%��5��������~���B���)z�x��s��b	�NMPm�F��A�B� 6�G2 �2.�x���zɁ(�(�=��L��גA)�P��'e�����`�Ka�s�`�K����_��(w�J�j+.�hN*in̉��& ?0ꆘ�p��QG�k�׌�L�H?:?���%M�~���ҞZ�M�����	SC&(��Y\��B���;�(/o�?m"hgl��)ؚN21�����@�'������x�擒���A~���0��'�8SH%�4�j3���F��<�G���-x���0y�jsa�L9�U,�Y3��������e��WuoɵE���A嫻�7��ݷ��pc)��܊'��9��w��>4�����¨���T�7�_dtS�P�"&r����.Uǟ5����m�V^��� �1����ߋ��� K��[p ����� �A���>�K�$�+���1c�@�/�'�]�j,S0����G��w:�*+�5'Ĺ��H#� ��+0�)�/[���EM�-�x���hι���y��#�t� g`�bmj�
�c:<���E��#T�L�n��9r���!!��Tk��^���w�/�i����@��M�d��.�����9v}O�E�6��H�f�I'%����*sqbn��i����`�0��'�?��4�w����;����/�[��>}��̀8\'�G�z�PS9|#�*�#�o�W�~O�	��U����M��հ��6�����7贂�7���|�R�#�]�8s��F���t�ܾ�04Sa��+�T/�B.j���󇦍5���ɋ�H�?ё��CX�JǜQBfa&�jȺh�ޝ?qG�⵻8���PX�x↳m��)Z���7�-��P��-`�U�|j	W����s���!;(�U����E@�ka��`|P:���a�ہ�ƀ�-K�:��nǜް;�/�@dR@�����HbB�O����E�+1�·�S,��I�<���N���h�����v��gg�N%�t&��5�Hà��oK�1�@��7*�-��D��z�fĳ�v��*]�@�R%B!��Bh,f/��8�vŕ?"D8}�yaQ��q����y����L�-��8��6�,�zօ��S��pR(Q�<�$H
_nYA^(�bh�>���w�mơ����Х��Y�[t|X��׳{5���=~�;�|�߄O���fO�[���Vfaw���˛P��v�\���g?SJ��XC���� {=׹Iy ��J�ee����R�QZc����q:���xl���=2�*w�ȫ�)]��8o����+� �n
Y2r�¬*b*��v�r4rc,O��+���x����t�'e��`��C8.��t�4�$�㢓rb�>#���\Z����n�>Vjd���5ʀ�NN���E�|�؇2ٛ� �1K�9��'w����4��+��9�0��XNE��h��^�j\�3��hWz-I��&�|8�~`��4�����]-0�vh���@��߸vO�Xw���I.�t�+��D�^�������4^�@>S����<)( s�A��,&��à/FA�ӏtx���t����UW�s�`��R���=쫀�b>��60�����<�ԭ�5mQ<�j�V������m(�c��j(���8�N�����@�m�L��yOń%�܆��p��ⶠ�<+K�M�����%MB��Z��$�u	'���A �y��N<I�O ���K�|m���Ȼ�*q��uI��,'�Z;���9��]ʈ�J�����[uSw(0�_�6Z�`�,p3�i�:��hP6q����9�S�L�y�]�" ݜ�GA*��{#`�e��9!VZx�jLl�;����rĒM���V��כE���	M3�lw��c��"�(�U�J<�b�$Dְ?d�y��Ûsa��?$�iQ�*X➮����8�j�c�<g��WYv���a�ғɁJ��E��J-C�@l�y�R��`aP��P)C���+w�	������ ��H��(��蹍�̦l��
.�2D缣F�0�Gdoo0��7���[������I�~���*�EahG<���)i��WΖ}��wČ�x�z�7��7�0�n*&�ԅ|e��b�OQ�]�J�!}2�щK:FOB��0~�]�'�Փ�ȅ����SE�|v��k��O�z���1��6?	^����"�Z;�>�z�T3�9'O��o��6vt�]�O.XX叀0'� '�|��p~W�r���E�5�4�ԩ"�!J-�'�Z
N�4����L9���f~���V�x�$��邀�n�s�E+��eZ��p��{�l�+���cW�m���U�>����Jo�2~4?��2�����\�Ӵ��{�?n�įԿ,T��!n�sã޷��×�(���h?���|*Օ��qÒ�*&IO� ��Ͷ9����	���Z$��gk$�#�g���j�a�2eK�߀"��5�,+��3ӽ���y^�?ͺ�Wi��_��BYבֿ+���F��?@�����f<�o\���[q�K���	��e7�v:��<��1�Tp�C�yM$���M�DZ�_�r>��g*$/�z�{�.�*ڋ�E��i�oȚ�ID�mF:�%5�@�7����:WG�%k��+��ʍ2@�{����"a�\�5YЯ	���U����m�wg��ɱ��?�JmĽ0�9L^]�,���sc�wX�w�q�O�~1��S�^qV�UvL��	�5�E#TOq�3��H��m��\`T5���K�Kd䁫�p:�v�L��6�S��S�!� X�|��P�ɫ�[(���'��z���H���]"�"�~��\��Fiș�yå�.��[QF��޲��ɣ&�f�ӹj�[�D��4Cߑ��� ���o +��w��q;�"���2	�$��)�x@� nO�*�"���&-΅;�D�q-#�\k[� ǔ���ݧ�i١�7��"�q��3�����[;����ۧ�ɻ�`����l�$����Ʀl�j�A)���|�L�#v�7��� V�t��Z���6s+�޷�8坽�X�vޖ�S�沬��P7�<*�Ütf�bX��6��D��sj��f��?ͳ&p��u�=�L��q��]��A�
#�ޒQJmt#-���`9}���+V	7���YT��wֲ��O*�C��;~�ϡ/��e�9�װ�L�Xi����%%JQM`��5�Mx���0ůx����(��4����HAU�F:��v:��,+ąɨ����4�f�Q�.\=�^�P��a60O���)�'���G��=��->�HՖ�u�Sz#�ݡ
\�zꞿ�̝5.�S�U:S�)M�>�c�G q`'+=��gY�)�k�a��LZu:"� �9h���{��|���)�ߦ��Jg�t��K�!����\w���|�-��r�l���?E�%���L�eF��&��B��J(5s��yɪݦ[����."�M�&��}2����\��S�zC�|���W�_;-i�#I6 b�Ȼȣ۾���Y����ڽt��S�DO�!��7�3���av\�����t�`��*4�=�	'(l��Xm�\]*Nڸ�N��&��dDXh�}^���>i$ke^�ً���Gu� ���C��b{�+�zqD�~{�O�0M"��W\-U�z\�e��f�����X>s���5��S�J�
��Jr�Q�+^�0�&W߉�Ļ�]�œ~�W��8YS�M#�����X��Wf~����Wk�q��pʯ��m��Jg�<�KSXz@_nn)Sg��)V����K&@āń�e��kU��v�KHa��j"$�������P���B+���k�椴�����D�2,���a�A�t\�4��!fN�$а����P�&*'�!�[^�9�|gӻ��mŋ����	I*������_�`dL�/���k����h"�I�y6(W���E�Is� tǹ�O��6��r5��N�<���9�U$8<�%l��t X���]���U�B��K�P{���1�g�9 �9)������([Q�=�Al^���c�*=���o&��������ӛ.m6	}��c�h�t�*e���P�^�ւ}���]�Q��aF���AIc�2⁽˦�k���PW]���fK�Y�e��x���1v���'ɐ�1i��;9z#>�	�UъDN�C���ar�ع!r�Z�"K=7���a �Zt6�?1D�mLW'y�xN�(79�������ҷ����X��ܛ����޽��P�e�Ǝʁ�C���u	��{�x_�a+sDts��DF�4fX��+����~E4��qc�wg�\�y����6�i
�^�|+ �:��E�O�,h&2O:?!�P��X��ЮL��*d�SP�=��=6�Y<��qXy+�u�Du�F$=�6Z���% =�~/�CZ��K�cIx�TJ�N��0�����>�qh\�~�� J���KG�����M��X/��.�����נ1ra��M)M����j�f;�#��8,�]��G�����	zn����	Xx�Z��l�Ȍ2GƎe����G�u䤹k�U���:����m��"�2.:���c�%N����x�GP0��b����V��S�"��Oz}��j����tK��n����"��U��~K`�D�C��n�e(��Xe�H��1�G���J;�7աWBy-J	���i�m�l�����, t�ؚ��ߑ��sW�s�f��V�X��pA'��	x ��p��1g��P�:e�gY��nщx��CЬc/� ��j��*���;��?3�2.#Ҩ�x����:���_��	2�k��6�r��2O$�f��˶����r�9���m>������[H;j�tS����a�!Ħ�,��F�!�ص��ֲ�ߗ��-?�� 1��T8,� ��g+�K��:��P���IL_���(�b��7(��Պ�����s���G+��9K<}��	n�|U����¢j�H��ˏ�S5���Po��р�_�ƛH�L�c�=��h�|��E:wIi�+f�I�zݱc'�#~Dv[�&�*�!e��1�V�J���C�f�*z.�YI�8v��o�-�Ρg�Ǯj�"~~s�&W�b��sܪF���aa[�����~9`\��bCO�ӷ��}@�% ��pJ�U�Tk_���[�v�^���0#�)g���T�u[I'��`��$��#|*�����r�&��f�ߠ�yCnN�¥7����"}��,�cd�.J�t�	���v�l�۾��q{� l6��
�\��r��:/G��3?&7��{��X�4���Hj�+�-<��BA$�>����oF	# "U��=��RCLH) �p"F���%��6�B|��V�\�9$S݉|ю>�����Б4X��I����^Kcu���4���T~?j�����i{eĬ��Y�c���F�!�{|�����X�V�������س��]"K��_H��ͫ���n��I7r]l�H(6���0�i��qg ;+F�Ai�����������Np!���M�xg%1&�*�2E��מM-L��=-R�zo�3%�Y������ޝ��|sݛ��I�_8[MI�����Aw�oF]�4�ڴ����xז�,�k6�\����GՑ�pbxf�������`���ؕ��#�Y3�r�&�ı�7*�i{%-?vd�}}���)�a��q�&����6���a�����k�ɒ��q`6@� ��L�X��ő�W���j��e�w�H��J�.U�R���c�z�w1��x��b�2mU
NXr7!�Ƶ��UZ�<���J�$9���~6 ���N=����l�����<�ʘ��&lYW��o�p����B�(�EYB�h��hO��V�o��i|�&gRS���moH���Rm΄&�6I��qI.+k�)��χ>pA$�@o��ϼ�1c2��|}v���JwJe߂K�	����ڻ7�׵v<�>���WJ��'��.:��F<o�����A��8HF����vS��E�t'�Sɶl�<��r�Śx7ǽ"��Fd٧n�w���y�MD�k������}wdF�x;:^�k��e&�	M�d�\�Y��`m�����]{P+�1�+PSi�c���7
ӥ�_t-pzm����!���7����|����H�WS�(���Q������!C��Pj��5ȕ���A�G�i��՚�����R��5S�lV���؀�~d���ԁ�eN9���WL�
#ȗRq�����r���R��f����s<~ōp�B�Lie<��ѷ�#�=	ĸ]r����B�"���\y�4�e�.�b|t���Xg�0o�R�Y�D�����X,<ͲLC7� d���V9,v�@$ʺ�!wW],~�_�7����|͕��9m��5�KE��d�7�'�jl��P۲�NS�*0����=�XO�xG��>ԁΖ�qΏGr7Rv��y5�`�΄��6�#��6��C�cg:4C]�������h#�	vD���ӎ�A���1[>�"��VxTU�����+�y�o�79qP�����b�h� ���1�"�h�&䲀d<^-��$|��/��#�>`\����6xmW60P
&z�5����K�Ό���ݝr���Wk#�;�r��ڝ�n�q�on��vkbl��A��e����Yn������[�h��M�Oh A�c���-�ڍ0hP����K\�완�`�`�`ۆ�4���"@q��U&/D]T-�yl�
ES�gv"���I�zi�����- ��S�S,=n�vW3"g���6-qw��ϣ@�+k�N��Kmc�G��L 	.~Ψ��~��\glpt#(��1�.�Ҧ���i�Y���\��.a:�׮��G�-y��g����ʹ����������̽�G��I��R����Z%�QC���'e�S��0eB!�9�Z�vi34;���-�!�݈�-��VV�Lzw���F��a����=��Ԉz������1)Au��@����g�z;�n�����	b�/ Z*	�B�'$�c��1'GH|�M#0P>k�����������K��O5I���tAYJS�s����8~��Y%]8M��̤aM&#$���=D$9�&�G~Q�NF�:�=rZm{45��E3��qk��\��ZAŤ��� �X���?[]1=�<�y�[�U���We�'YĮ�?7݄��'���{=A�Iɳ׷��l�Ps�s�lB�)�ȋ��
-�ȌP���qʥ�ϭ0]���[�#ulA�I��n����ZB�l�Mn��J�R��Ww"�uyf n}�����Ux�����ql�H�o��Q4�B�x��[,�*l�N�12��~�����t��N/����l����yE���-�����RJ:��۹G�����
����O=M�S�ܶ�ݺ���uS76s(�8���@s��Wj��#(�:��iEQ�,��~�a��w=�F���kt�+���$��ʩ�rцJmkuu�iL`U��Xu����i&������s�o'%�;c��3|+�Sa',ug�繑���[�s�@���a�;lA����I���I"�2.�&Z�q{�"��3��-��8�X�n�%R�ԫ��M���v86b�<1Ț7����Gf����L����(*�������Ⰲ�/8j�M�k�-�W�p��R�R�g�������T���c���8oB�>z���}��7A)��~�"�5Y"�&͹���nU=����Li�zS��d�+D�{��� 10�~\2�Dn�C���1˔ͷk��{��L}o�K#�� ����Œr&`�Ź��x�j�"��1�*z����@i�h�|M9~ E#����.��Y�#}�蒬L&�Լ�M�#.21�9�Y���l�%i/�Z�LR��(�3�;�HI�ql%�)��u◌��
>\��dC�
�	��iv*c�ӥL�K3㘬�ԬFh���#Ɏ�C�O��AZ;��D����#B�˙��2���	�����ħHpVs����O}��_�m��f'�W�56G�	��������Q�t�gwy��nu���5� L�Z��ڤ�[�`[_1i m�rp�y���ήL4���̿����Xo7�U�ů���;�����$�IZ���?��"Kt�l�����!���䢾T�Ƿ|c�Q��A ��S{(	y��[�0�P�l�("��|k���d�5�A����M����t�j�a{� :�_XZ����pLh�'=���.�v���j���3?�&��I�m>��/�o[9̫%�	���L�&h��X�ӡC��"���»-�?Eںpfl������e���fT�T^����@��)�[��%�M��Y5��8W��#K���	�r{�ޛn0���ʹ�?o6R@ ����y�v�t�S���S9������Z��鐶�A��gNH���?�cB��$Z�u�R-.ͬhc�.SL�UA�{�-evBA�5_�석�}b��d[LL_��q��q�`��Sj�}�>��i��
��R�U�f�I|�0_��������B.<��4�y��m4���n�������ob/����"S�7K��0E"��(Y5�hn4c�M�IQNL��eN}��2 l�ޝ0��/��QvP�-m���7n"�����g���v��oS��qu�޸�wo�7td��Ȕ�*(��u�:-�����Us�y&�}�����J�s
*��Q�ڞl.r�uښ�����r�Hm��͏h���@>p��h��IM����Q�x/L��,���F,�)eVK��|!�k���5�)�w8a泷�Ɂ��?���]�$/E_�Ѕ��
D ��\ ���t�|V�����F�]Iڪޅ19"*@���Qkə?A�p����i��B0��;��c�9$��gRg��4��kT6y�'9���SXծ[ϖц|������B[;d͠���^��4��<U� +�0���@N����r�g�62�ç��I�v;��LU�������h�4�����z 7��"��{E����-���+������	�r�<S�=�p��P���
��+���\�G�y��ܙ��N�[`�}�(J��bS����B6q3��lc�/0�!!�݌��΀��K�A���[%7I��� ޻6M�=|���2w�n�Rvӵ��`�*��<x�v>U �;Zʦ�=%�^9_����wT���967����*�!��5 <].,�����I�^�h5�!�/+�:Ymc{���_$b��m��ϫ�]�z��d�y�g?Mu����5:��&�Ӓ��e�]
���'��"3&S�!�s�m�O�#b&uNG-5����zH�<��"Y�T�~pГ�$�e��{�X� ���0���w�hcK�5;$S��KZU���M��۸�����=���Y�S�ȿ�U�`�y,�
��/���Sw>=C��	)���Fy��%e�D�
�Q�O�7~m7XޕJ=_��6�.G�9����x?���6�۸C��L��}�(��^�U�!~��T�3L����+��� �Q�2wLx.�
9|ZE���:�$l
6���=��(�� �)k��;`s2���q�t��NM���d8���ড়�]��鵁\�4˅�웛_�%�-�埕|�02O�2G�r1��y��s�'Ǹe�[����h.O,w�@�؞��ߖF���}䃇9h�G��_��MG��;X�}�}KW@��5`Wq.ᠬ�y����|��QN�7�6�_d�B ҋm��u���$�{��!���؁��D���zH5hLI����D]���j�"q��(���$����3q���8��~=�͕m2�(F�XzB������ĠQ����nǞ�B")�h�o�ʹ4�1a��%���ٔ0���w��H�9�ϕFnJݤ9����k"�^�h�aYh@���y��;�O&�����SG^�"����R�qR���7�����%kE�X9���?D���A��9�� )�6�-}&v�'������dG#���Hd���t�Zl<���S�Q�eo�uжF.�]�"`���&A�|�cO�b����6��<�O���D���"�e�v�K8���4K�,N"�\ad���|��*�*�~�#�pU�߹��u�69�u[,�T���S�=+7"�.0PdjH��A�b��8�m\�wQ���M[n�t�߳¤b�Q69�f�Qt�V�!@[
T���IG�F����q�֔Q�Ǻ�j޽\�����|~����be>��n��Q�Z�#�$�:�x��gq4xG��
�����(WH�� �%Z�1�����G�/B����\��Zx:5��K�Y}j����s���'v��O������2��]�i�S^��DWr�Cu���ۇ~X���4�w?�<�@�Ea��U?��F�����c��KP���0To��C��)"��T�#�O3�T�v��&���48���9����Й���Qݍ��ZǌiDi"���׌��+��k|k���ſ��Z{ik�u[������V4�,��HP?�Lg6�E�5^r���I%�>�,�����Y^�)�e�:]�G���lz�w�n9�(��ߞgW�(���4��1��I�m����f��N��G�,�����;�O�\���<��o����Tu��:��.�D%prp�R&~?����֟��2��s���31�S�#������phv�_Z�!�o,���62m$�^+����y�U��d7�&R�20)iٶ�;{R��bI
a�=�}=IYGG:.��O"&42
����8M�o([������+�N-A�l���Fr�fQ���+%���0�æ�>"��m�MR/3�-l��ý$/�Les*�+�j&�޺ߢ�,Vޱ"^�!c�1f���iH�X�_G/���8�)�hiT�c����Tt�k�B'j�b`w'�I�f܊'� ��|�T+����`qժ`ǻSn�_�o&��������?Ru��P@Zm�ڂ",�$��w�՘��e:�6[�yl% +��J���q�%`?Ui�aҤT�����K��5�%��B(��QA�O���<#���ʂ����5�����
m�W0;�o�?�	�H}"3�N� ��2�׳��.��0����9�U��#�vL�n��>��>l�{��Bu���h�r�J#W���ԁ�f%��1Fn�Y�<(n`����S�gyZ2�_�w?J���j�m�	7��[@��9h
�H�L���&�� �\Fuum'Zd�E�.��sd;���pt%u�>H������6��2 �R�q�6l�gڳ\��/�~-�Gd�M�O�}V����]�;��������
PD5��6g�`�]aO4�2 Q;V3gzx������	[9�G�_Mu�	��i��c�����b�O�:�*�'�BVz����V����"x�� CP�
��`�)P.�ֵ�t�qz�J� u�?<[	c�΃Q]���W]ã����PM��� 2Ɋ2�N���fD���~���ΰ��b͹����4���J�r/]JM�l��,��"Y�X��FJzCݖ�H?jc���������m�A���յԽ��ϣxuurϵ�V�Zә�*�G�|�	���V��;$��!�nxF���}��f' �y�I��м��f6��3�8�xD�QE�p���8P��H��N5��FM�
=%�O��;)��&MpQ̊�k��������T�|�����l�u�7Ik�c��_���Oeזj�&�Ի�3��ۙIYE�4�buȍd��XUQ���k�]+��'�X���%�ı���/A��{�LY�jl��I��I�}�p�	I���ǿ³Ly�e!Z��IP�b rpA\��M
�����0
�XJ�n�E�v�yT��&fnK#3t��{���!�n�Օ��������>f�A*�TA\M�r6��o�b'7ߍ�D�����pm𼦩$3�/Ȼ������'��\M�O(�s@��^������v�{�?��j�fi����,���ٽ�~�wZN��̉�m
h'o#�DO�#�������R[I��� eC��8��7¨�j
O����`OyI����O��7f�W	;��qX�Y�T��'���`b�M����B��7�R�7���Q�J>12&�QC��+8�}�0�VE&է�G6'
��k�����R#�7&��:�v��!�̳x��~�Ę~y#a���:аLV'���uT�{RĤ�j�ƙ����iG4�P�����F��FA��إ)��m�Q����qlŒ��h���P	d�Gyx�0q��MY�¶��2�0�u��
~Kq��@����h�so����H�hB{!RPv@?:[��<��ĭ�
��'�Th��U�줧�c���'f�}�ĸ�W^�!��p�u��m��x(CU���`0,���k�8[��r
��ڷ�Ƙ�|��(-�l�����Z���7��S��V0W�t#Vz6�u!�i�jt�ܾ�`Lr޲�)yq5W]r��zܰɼx}�F���w~�����zc�G萘b��1��5>G^�e��2�
��ш|��w�f1'��\�2v����n o:���*~OW;�A��C�cdX����y{Β<����Ǩ%Y��a�e(Ry�)a G�qu&��n�r�����ъĔ��=-�W��K�Ed�q>?6�\����R�Z��|.�Se���%������ �MA�T����'q8��x�)gۆ>����#�A\6fY�����>[_`T�U�� �z��&���f9L�1e�>6\�V�X9S{��QIS�6�x�*��x� i~���Id���I�	��B4c����ብ��\e�j6���psy���8$Ö.7�Q?�vD��?m5Nyc�&�����ul�I\�[Ot_�� #��ym��ԟ���Ì����99����Ώ�a��>r�BA!ԑHx�)�0��=Q����nzi$�e���#�1P���c�B�
Hj GJw�9����6���ڐ�1�38 .�9"�҄�����k�[��f����w���!P���?�D�F���aq*�M����� ����]���G��?Df�I2�,��]��1�&�������G±��������r�(كdn�j����q�(eG^�l�jv��8d͒���[|-D��'9�b�Ͱڤ4P-��u���V��[\�r���[m���@�}��8��S�Tk%jgp�x��X9z�������b4Ē�t%sc�����{P�X� ��~;$";-�W�Ƕ�>�U^%weQ�RC��[C�j�;���I�9��m0�߅-�dy*L-g~F�?V}��״p+~\�ǯf���I��7��V�Y���Ml�����z&��AV���X���qޓ'����b�_9��M�a��
��8�]���Ә-���lda��r���P���"@�s�H��M+�X�U{q^�_tbZ>X�G�&����r8��y� ��G$e�̨AFc�v&`*XP_*��X�e�F�8)J�U�'_GX�Vl/�(-J��kjSF��2��y�o�(��X^�YD�MF>l�|u�R7��E`�?ӑ����X��GH��X*�>��O�B/��s�I�{��2O�98%+G�Qڰ�֚�*���>��#2�J����qÏ\t�?#����n8��K�_�� �/�=+��Ϲ�'��3p���Ŕs���"]�Uھ�����^�خ*��3��=��ًV�x"��EHH;EoIu��~��O�_Z1�~����ĳ��U^"n�H L�7�O<�2r8z�N�"w�aLnM*���i^D^=�Q�"��bV��w�He�֕�2��&lj;aF����a��nt�t*u�3��j:��e��xmA|4��hN���%@��`Lx�XW�/�$�TD�E�+A��#�~e9zȼ� �`�:(�|x{��_� �P�lOy���R<�5�z�9{��ΐ30�f��	��/?�k}_��h�\c�M[qK��ˮ�`�ED�6Ͱm���8�Y��w�&U�}@�[�μ�ɕQ�Nk�Z���>��7�U������)��2"<��Tw�TX�I.|�nF��b�aQ=�P���7)Z��2<@�}�=��F��2�`LS$"i�����f0�����yRD�N�^ԝ�\���^�c�x��g0��(`׊���ߠ����.�L1��z�e�6��d�yu�m}�䉏�*�{l���d����'m�/�����U�J��r��ĝ/��+��5�S%�4I�q:st�N\~4�}�����+@���R��ct�&��w�y��`Kw�x2`�!�� ?W�)��A�u��G�YU ���}O�hi���Ֆw7('��`��;	RgH@�!��zv9��_<~f-8��:e��ͥCq%�}R�@�
�����l�=Y]'f�����r�K�.2̹L���|]nT;�p�$�>4՜���\4{�@��n@�
/&>��J�
�? �g������P':~x�B^G��5f��ob��D̽���w��f����._���������W����Տ�~��mO���TH!�,������6/�?�{�!�eS���Y?�~m^U`qͩ�&7��~3��Y�;���Jҽq��3�/D�y�l��q���M�I񨞐Z�m�k�����O�>�-��ؙr�G��Զ+ *��Y����Y��;2/��lao^w�ظ��~꛰4��(W����۝�5�Y���_QewӸ՝t܏B�1�R3N��|����l�&^�������tߓVL��,Nd�T�ѪX��Z��{�;�H��J�Al��,���(�`V�x���Ri�
,#{ː#�W���(��j'"�� ��T���'}u���)eG���J��.s��\^(��Z'�Nc2�4����ۺ�鼆��@���)2b��<�o�	A�BS��*t��=����~v��D��Oz(-cNm�����EN	H��h�e��D���~�/��l�ʟ��?�������љ��%��c��R}����扇 ��ܛ���t5;�)<��`�!���w*v�����p�'B4�dQ�)�fm���a�К��X��\����͙}̲��]�Afe�;n���+�~i�R�l/ڒCM���ʗY�����I�T���À$��Qk.�:� ��c�E�ǒ�s���H��kE�ł$6�G�`ߙ��9����ˁ1
fOy�	-f� 2�J��Zt?� ��^m��{h�֫��a�):�#�{2������0+�/�k!��=�/	��<�ra�4�����)V�ج�*K�b�񅀄N{�>Y��c�l�l�~�/��:5�ee,6�]2�A�ƖZ�gZ�L4�>�����/���\�Z|��)�]MnǙ�@�7�<P��_����[r���P���'��B�qhji'��r{Xl�2�rvz����X���r�J�4f��q#��Cu���*����y�Y�vG��_�tqO��Ɏ�ړs�q5��k��S�Q+��~0~����[2��Gǌ���4}g�5v�6¥������	����h�� �85��0���7�E�_��R�Z���)����1A�/�q�;)��3�`�'�uF�Y��\�Aʥ�ȾD���L:W"-�5��.�����������jS��ԄT�5�{
0�G&>�tzX���qJH����Qgi7��dvm�+ky��R�!$���kQg}�����J��@= �ꋔ��Wj��R���pl��""����m�7+nm:&<T�r���V�����D�_���>"�Y���+��X��罟~+�6}W�A+�u_-:�l��;���r<4��31��pI��1�=-Wk�}�w3>jc�y�EU��ݏ@��lA�+ �)�i�*�/������ײB�Z]�DwW�W���aA�M�+H��L���g�����Pc?���@w���M�z��%��n��e#e�՛5'��''�]|5�״��4��uYLK�j�qp�:��N�Q+kza�I�����w�D#�F���yI^_�%2DpZ�+DjA�� �6������ ��I����u-��9"c�T�9!-fu�a�,�qz���S��q��cv��:�!AQ���0s�I4HH<�����%�a#DB:~���{$��Q�����Q��}���������!���������.-"
�DN`W	�fdƾ��%\��N��#���#�`��~	�B�?��!7��C�r:СȎ;9)�]y*����{�h�։ǰ�����+�Ve �f�`Sз�Q1?^l���ߒ��� �����W![�4�m� ����=��lDƖt	�\�#�FN~8��i��o�R�ݮ��;]��4��%B_�m����$^)}��&_~�s������<!���1��}T�& �.���/M)Iő�Pb�A缓�I������`�Y<�R���5K[6�؊�4��-�'��\nB�z�(r����-�MOJO�d#o}xM���M������B6u
w�y��ޢ�T�`�k��v��O+[�y
������_�?��S��<|��8�*����5�G���ҿc�K\�S~D|�����Ǩ�n5b���e\�;gRl�A�܋P9ǟU��\��� ��n�w���ky�b_u����6�ɪ�.�����JO�	�&hF��S�aU(�7s�=�&�m��0��V���R\o�ކ��hߚ�-5��0z��
-�R����O���Cq�G�D�z���*'��i6n"8B�3W�6S�ꢧ�6)���ـ"b�X\�x1:,W�;x�9�ǐ��g.1C(sv��8�)���)�b9���2��#h����d*S.LAo���/������ W�*I�>M'#6�Z�w)��~٤�X�~��j�,+��R�[�.�a8g�?�u䴫� k�m��;*G%��6��9�́��C&b�����p���ݙ$Zo����#�i��&���(�%9���Y�q���1�Ls�Φ��I����Y��ҋBq�sc&���dƃ�p%����w����Q� � Z�ū@�<I��Ј�� ]���>t���wi�>æG���f�w�����J�j͕�и�@J�1�̯�tM�q���v7��v*ɏ���������M�eQZO8��'��a`��p{�Rd�?10w�t�mK�����0`��fa7�pz���'�$���ÀHJ�][��d�cz��pp%�#x�� eJ���y�f���?��B�b��P�ʙ��� y���|����-ܱ�+�"�	o���#gȄP"ք�Gə"���P^�x\�<|G0b��h��*���G�6 %�N��^&�%���K/�XL$��+]��#��{-���_Y��OU/�_�YW>ām��Z|c��跾�P}nJSuq�������)��]P?~dV�F䝟�\s�����$�^���$�%����R9.��i���|Yŵ�8m��(�u��m�� �W�;*4g�Y�t��g֮��ػ�b�� ~\B��E�^�.w$?6X�ߊ�ϼ�r4p�d�Z#<�Z��D^�g�+g�p3����\𖏌H���|k�=iVV�	����Qv#����,�>Y�׿/M��эK�as'\S	�/-�8jA1��k*���>%�w�������)����p��G������c�d)yoI���#2~�T?*�A]Q�tB�Ll�jfE(���/;1?��x�4�dw�o���J��d�Q$�sNfKp��]Bo7���i�:-&_�Dc�%L��"�eYO+�H��#���>y�yi�()���l�,0^���'�Ӭx
�'~�Მ'I�sù���!ha\2<��V�h��a�� *�1�'#|���o�L�Ω.ቿȮ·�p�����T7��Lo��k���T���W�Q�G�AL�~�;y4䭎Wb�4������v��#��Ze��\&	c���*��rV�z��?Ɔ��.��%�����G��03��V�H:T�h���K��A�eCu�^x��nx����I�bK�9`��`"�rr�\f�Bl;[�5*�@I���ښ��^PH���ʹKu��V������A��������d���Y���t>���z��D�cu�Jvͭ�?�]'�_ZD�R�.�Ot����b�L0#�af����6����e�4~a&�,��.T�K�lDPkK�f�IoW�y�r#u�2��5}c�π�-���65V�EJ�Ғ��w�mD!8���4��Q�+�?��8���^�uAC���L��.��c@�p
�BU
�>���ar)�����.u�׾_f���̩q�M��vw��W`���A,�)����X����B�d��Z�n��������U�xy�Mkr���FYWX�m�A�Ų�S�q�r�k6� hq�U��A^O�,�����L�y�м��
^=`��p��%\���ha��?��)-�K�l��Q}�uc�{�iY��z�L���_�(kv��3 ґ5W2���o�[��)n$� @[X���T����X�[�%*��0�'J|*�́�|މ"�Pv}['������o�_kT5D�+i���I;8��Z���[��}э�e��AH��������3�<��W�Hz-�j��~��ц@X����=����&�&&�ⱦT�DAA��X���`�z,��=R�G�h^�3�?�L ��:��m>E\M�P�R�=�2�ƃ��H�s��a[`L�g6����Q����$����&� ��E3:N�IO-mz��[�lQ���0�M&O��A�kx#6���'h��DM��Y�EO�'H`��t��7���ζEb�)�>�ϮC����Z��e��Ԝ��]��k�,t}�4v�[#7�}����"�w]�ͮs\���CM�e:�Ӡq���������O^�]��}s�R�
�&�N\��նӁ "�\�}�wU"i�<��=���	��s��Bz�����~��)̖^_�k/2�����Iڲ�Z��
S�@y
<FS΋���C\�6Y-��pb�������t��_��H�a�@B��k�D�S���5ˀ�j�$m�J�^c�)2KD�qb�qpZV�#�s]�
��ZEUq��D��'^��V�����Ҧ�k&8�˝P�����������a�N2my7�KO��r���`$'����nɚ�"�����2a��lf�vrtn �S_D˾�_�,�&�bz����f%O���
w�
 ��R�Ck}�	���?�T�2,��g'`�L�w})��<�ѻ���PIT؏���a��jI~Ә��3+[�����b=��%{�1�*�ujR���x�n�{䙘M�8U@�d+�Yd+��W%
��(,JQ,��18���te�',�dH�I4ȏ�+��Y��K���_�1��4�����({jP;��6�D���R�ڴ�T��ev���]}���E�^?��9�YG�Kz��Q��|4��<�69�~t{r�&�g}{��sI�������Yt� �NOڋJ4K*K�x�Æ�;^v���@
��|�!T����������T�!=%�,e߃�`�
��dZRv������|��|�ְYO5ZV��s�/y�>5ӣ��ei��sy@l;�����gA^ڏ�� ��Q��ߏ�r�s�$��SB���'�����WYbb+�'�tնʪ��&��#�B ^�>�o���0@�����h�d�Ҙ��bPdv��h�.L�aT��``h�b��ږ��L�.�ڒO�k{���I�Q�v�`O3����J�g>�s]�#y��v��Y�#9G�8�g����N�(^��d�Q��j��{e���x]��� 
6�v�=�k��#�ة�(+l=d�(\^�㳙�����A{J)9��u~�s�S�-;T�����"*�UXA?4�������s��π��D��6>i���T��)��$��V��}���V�VsP=J��Fw!��ٚ�[�?�g%p�#�t�"`�G����X�͸l>�-�{�ʟ#���H0ôDoG����ן��*�ugg�5$�0�9�γ��Dt�*K��X�����}#��\N-:
���*R�����-iY��k�H�p�9�&#;5��{.�_�@*<�Hd����PFۏ'Yy�B��u��r�W�^���0��/�6���k=O�d`�Ԯ��$KB���c+�e��F�Ȃ�l��E�VDF������C��`����<��j��]�?�d�@��`}�o�f���9.�f� ����S�>MX�أPW��WX�d���A%C�7�N2��?��~zYM(2���������E+����p��8��$z|��cCor����-xz������ƈX��dt�Yk%M)ͯ���*h����7��ш�&�Ycz���(�r�"WL�^H�X�m���}�#�z�pS��C=��@��q�f���ήޒ��?��#��g6�KJ�$��� E�qVs٤#pyXlY���Z%���rF-v� �b�I5J�.����t1䫖����'qE��7ާA��c����S�c��-x�G�EB	g��o��(�2%Qq�֞3m7M4���U�Mہ_�r�&)��8Ҹ�;�M�H����%O����C2�3�5[�<(�	bęק��E�=܈��K`��	R��M=~���|Pv��*H$�_i���$�0�y�s��7����9=�&Q���� �U0Z�v�g���*�$\��o|��T�u��ꗧ�E�]�G�k�F� �9��|[���sR��f:����OG>G,O1��#	�~�bV��������2$�5��+t�Q_z���؉0�Ws������X#���������/@R_4�����>>��q�1�U���3��H���[��Thٹ����
Nы��� )XD�%�Ŕ��������U��eD�+�Ք6�GC`�}}02}1m��g>����F,R�W�5���z0��L�/�k���":ܹ��<u�1�<��t�Z�ƫ>j��������na��ӄ\anB�� D%�5�Uv�)����':z�8�r���b�BK���	7n4ۈ!dDY|���U3�ݲ�Z���n�M�?��WB��t*�ă��G��$T�&�R�$�L��R���#0���(�]u�݈���-<{�V�}���e'sL�c��Z�x2�c�9��=j�Z���21?Y�K[m
Z���Q�$GؖU����P��\K�d����;���\	�	>�"��L'װha项�ס�9���\x�1t@��_)ϋz�l��9���kg�k��x��~1�Bw�zJ�λ����L�������?�Xt�}H/��a���P�ЋR���dIoGH_�d�!?e����"KQtJ	4Effx�:�oŅ[9�Q�?� � ��8�X��!�xl�M�ZE�֘Sx�Z���P1/:f@; sGԥI��9U��Sq�e��8D���m䘨��g�O��B���KP8_X$��Z� _S�Du�'Ѭ;O�;�Hݻ�������+p�Zdl��Y!�����s�Xa����G�CII��?Lstlr�	�vb�m v�.������M�NLD��Ѧ\r?�N�E_(zY�/3ЫT����8��9��r�T�+�x�1���1
k�퓡Q!g	���'v[���ŊY)e8���-�w �J����h�\_uA<o�W�u"lxu~�	1M��O��4/��������4R���5�#�Ξ�;�9��()Ք@�P%pwi��=ih��r��^�+��ޙ��t�6U5�������DZ��@�޼��=�46����ғ<�4?~�טWǲ�؝l��N�`�5�R4F��H��ۅ��?|"Q���&�|q��~��O�t�6�ܲ�/�2�����	%SK9Vw(z�?�k�R�1���ؖK]�� Jz-��&��,�ĺԪ�l�] ���	���1���k�g�r����Ѣ�+���W/�(A�)_<e�pA[DS�>:>5Ni'n�"tE�锼���0r;������>�K����1~�|/���G����V�Cr�c�R��7�:y�E���K�Ĳ1L�Fk�wO���N2��1Y��z�W���1�1?N'2q�E�J�K_��d�QhW�1\e��c�9nϫx����R�������#4L��,����e�7&����؆��óKOi�A<4!i]y8q����'��0�M�`ſ�ۏ$&;"�|vgȩ&5�݀�>U�~���D~f(׸�F���`c�c1��>{��s{DM����Ro|	�ߒ.�v�@���aJb�U�GUlC����坈�|ۂ�^9b���uHJ��#�Ei�����a�9�y�),����R&8qoke��F�pw=��=C�LOk]�J@�}S��u��0}*^���XXK�C�cb$��J�F�\[2%pC�J+���N]�!�l5)��O�t��Md�1�bfZP16���?����b4���
��Q!�>�vS���8�mlA*�f��� �j����.�#����|�i�X���܍R�������2G�		f`��綯��ƮO���(�e��Vj�4bc�{}����2̪�4���KuN��$�����|��4�;::�}iW�Q�X����J�WWz�?]�]>ˈ��������#�&��;5i3����x�ƴy���xi%�����0!�o��3���a�d֥���Ȓ)���D ?���9��85uiR�ݸ}s�rnL> �e����<c]P2���`�*�9�6s�	��$����%ʼg>��2}BuD��~-��Ix�2��!P`���e�+��+<XsGV���2Uޞ���O�j���؜�5����e�TX�q��6󔓰���}ܪ�{8He�lO����L#����E?'�����};�S�Ӝ�������-5����0���]شTZ:�ᐱ�X9�.��L@0}�Q+�����&�ɍ><�鹊_W�٠W������M��ok1�ꛛ
4F~�G�K`�dd����m�� G9�Dq�&�����;�-��V����\���g7����b�XD��,���������X`�����J�T����� �5װ3�M�pJ�*��r|/�lM䥨��q�Cԇ42(�=�S/ ���K��Wf8��N�*�sخz��W^<g�ß�v�-0�����������w|�嵢#Ø0&��b'0�8Ŵ\��͎S�l�oaex����K��� �zlnW�2���f;~M�z��IH�=��I5ץ�|�/��=-���Jٳ{��N�ߧ�p���͗��"��r��T}�nBas���cG��B�oK��͡ğ��W������F�w9M����|��RxA�Dp)�[j`J"Q��s?upI��#��ℓ�d�o��"�X����I��	�t���A���j�1�� �� �ٕ�E�$	N�������#㡞�̚L�?-���1k}���B}����Q��|���I���x�<�$z'N�X��G��fEJ������(/1K@t�0� BN*ث��x9�dG�� ��I��Sx2��7#.�k�@R"�cA���Yo��U��z���v���	��.�`=�Y��
D�-Uq���y^pO�|���?����pϜD��I����2���$���1�M�	����5n��j��O2r0�΋, ��}���r*�k�pB۸�]�<
P��_;5�82#���m#���KU�'�4��'|oZ�"R��'�rZm�#�W�M�(�km��khYLc�l��]�>�xC1�Y$]�*�ss:u�uH�N����R;���&Xz|�qsdS缼��UF���(��z+T_�b-����H�M��w�+����U:=��Īl��'2����O�|�R��mx��y?�ˑ�D��8|���r~%a�^v@C�����<��t���X<"p�B��5�ϔ�Y��&�cyD5�U��fy��>�+����Z�I#/��b�d�f���H��߹��}Z@�;����|�&���M��v}r�RT�Ԟ�L�JA4���-k�!=�m����a�t�DI���k� ��^q���at*���D��z]�\Ҳ�7l�*c�{�}v��D}M�煐�f@�&�v}�����|X���Ft���[!�ʈzh&����/�'��#ۺ�1�9Z@�Ѩo�S8���}�/ڕ�9S�Ujj���OL��3T�}ٮ��ơoM,�"�e�}�·iG��א�Ķ��F�� &��^��cXnuy8����o>G�;������`�bQ��ٙ+'"a��<�r�8�B�ѱ��"�UZ�M+��u7p(�H��%}���A1�t��x�dLW�WT.�}�͒�*L��� �����*�9`�V*�m_1����}tu���R��z:�?RPk��;֖�R� vm�+s91cbx�(!TQ�O��Leّ`�|#܉<�4��i�g��vHH$卥4�X(�>���b�[�Z��Dj�/w�Js�~8��J{���f
Js�N)t맺�����~L�����[�{�O��7^��>>Mqz9��Ԛs"�	���7�.�Űt��W� NO	��S�/ݺbK�s�!���LX���MAO�W�$od`�Uܻ�Wy���l���k�֢=��ʘ���&��%lq ���P ��	�Fd=յD<����-`����x�nB����¸��5�!
����0^i����\6"<H�&@3t!�/%����i���԰}�ú�C��s��I��+��PI�m1m�bB/Z�b�< =�������Rx��{	�,Q�&�|�8oAķ{��M��$N��g��)��'�͌�����}��_ܐ�e�=ӣ����2%!\;�0x�Q� =�YN�����A�E`r�uO?:!��Uw;IW�����Z�;k/%���d�_�$J�M������b�sCL��4ŮA�yV0��z��"c}�?�w
#��l����0z�f�:���gX�8�u�(���Ӹ6P�n��
��Z��̨A�W�f�P��gx��ھ$S�f�#�~tQc�5�S�`-%���L'
j�8�N������6/ŷVͭ6n�L��=>�F`�k1i]����SK�	�iЄҢ� m?����A�� ��[�jY�=W��9�'��Ԍ���۫�
���'Y�
�C�*�9Y��/ %4ۣ���|1�B�T������(^��E1K��0|�����w�x�<���%y
�.��ώ|�GH�?A��t�#����,$��C��^H��)u�],8��3����+�6�rP�m䜢��>+x���*�񁌯������WH�)�ʫ��h�q�q<����,�2��t�0�$b}��cG�/�wp�q��+HA�.����L5.��K*�G�*k���ݡ�{U|o�՞�כJC���\|�Sy�Ճ����w{V�["������{��M�7���E�&�g`��g;N����Z��	Y0��A
� y��'WMK� �I�?�Xr��ֳPކlp��|~N�2h���Vml۫H;M�vv������"�y�BQ�?Ȓq�q��S��Qƾ��lpD�*HV�#�ʌ����+6��75��� ��U�tU荕�Nr�M����`�]��;�}��Hѿ��2k�}��$B�cq}k��*�r�.�H�IjP��<��&�����N�~7��Lc�DE�9��`����K?�����V�Q���<���7�gz(~�4��xʊW*iڔ�6�m$%�L>,�P�v7wd��gޕa!�z��m%f����L�iY�<}m݆oJXp~�Ʉs��I�	Vϛ���Y��\Fխ��V�%��}?�~��z�Ũh/9Տ�Yj���.D����2�EM��0�IF�G�SC����m@@#�^7T��;�BO�aJ��C�U��u�S����2��i�n�ٞ�Pҡ�o��.��MM4�G>�Z;Z�)��Q��~�OQ�Gԛ>V�R���6F���]���� p�]������Aї�4���>�͔�U:7޷M�й2Rݼu�*�G0�6���%���`�|�ĝ��	'���np�ʜ�5܄%Q �64|$ư���P,��?l�\�8��uƎ���'��-�6��*/��jB&~����:�[E��Q��*�����cMm��������� �te�W�
�(���9{��:���Q$���n�(���}�� 7ciy�y+�n�����L �EH'���lL��ہV��ac��Ǜ�	S�����A3s�{p	.4YY���@;����h�� �
`vC��/3D4d���i����kKc�yԮ��$R'�L�)��@e��2O"������GDy�:�p��bs^�િ/��<Y���Y�䀹���F��G2��;6���0̐'!e����-H���|� s(JF�ES���e#�˙�>[����%E���cG�����yB'_�Ҹ'$�
�_��}A��6�XYV������촘��me�zď 
�	�H @���9��)��B�e���u11$'�U��[���Q���(Id�hO� C�x�p�%����s2D��^9�'lF�)R,�s�����AW�>Vv�@6~�܇��e�t�����u5g�޵5/|8��m[ϊ��!ۉ�f��cR7? �^6�_45U�@�]FX�jK"���O<8"W�����NR@`�jk_�0���u��t_E7�v��w�TĶ�u��-�,&�n����液{��>��W  �����Y���R'2�+�2:�ⷉPpHZ=���0R!5@��~/�ɻ.Q���n(�7ɗ6R����f�0���_��T�F
L��,��2 �[�q��GCS��Q�x`�R�f������D���Lv�1����Kl�dG��B9`b��p͚D�L��!.�n�|�tt'1rώf�~����vR�(9�a�� �1���\M{{��J/����w9�'��K�\�o�����c}����a��[ �����i�ih�9�>���G|��X��i�THF�:w�
ذ�yWj�ǆ`�,祠�^���gB�4S�kЮ+�p>�HLI� ]��RĚ[@J��d���ɥ��E\����x�C�m>��?���³���ox�����8Q])�g����m��s��ŗi*�-R�%`��� X�g'����g	�b���R��S>�"�x"Ɗ^	֔[S��W	oD��]��'5���ii�h������ⵃĹ#����:�a�4�(�瑙Ϭ]�n/�a�,3���xq8E�7�F���wNw��7�);���>`Ҙ��x�$�����$�y�RZg�Y�S+���zk"�v �|���:����|?��N6�%v�󄗩�*W�ov�R��m��^��b�z���J�3Gh���`�MȲT�����fT+���⺩�P�WΗJ��d`aC�3�sK|Mc��i�EH�sm��ז��'��+�����YV����Qp`3�5G2*���SG]T��*!��̞f�@�Є�v��Ly���J�t�a����y!Zkʧ�:�3T���_�jT{��v�ڝ8`b"7Cu���L��L�����H]�͏2G��k5���h��䫑V�����dFȗP��o��27M��E)Dw�?���h5�N��}h��O��XqZ�M�L��گ�t�h���x$��T�|��Ż���>c���M�ȎF����|�+��n�
��j���F��w���?w_}_�Q�5�� ly�����i\��/L!��=�1Jd�A�Ҵl�s��T�R�Tb������hJ����=ߒp7F*Ն$���Ϋ�}�Q���艘'�kCk}�z�k�;U*ٔ� �g3ĕA�Cb;�If<.0�y
�";:�P�2˅X�q��/�<?SܨF�2�k�{����-\1���#s]�"`s��@��x���Y��}-���&9!�v�4𳻛���p�i�L<C;t�
�Nm��E1�T/W_"d�t�ٟ�^�4N��M��U�7�ȑh�e�yW�=Ί2ɘ>���U"�.A�iw��^5�=IS�nD����9��"6��Z�FT��/�a����s���c�s����"��(@���tBj"�М�5���Y����n�|@�����>�� ����=�0���G'�=�|���vQ����f���݄qj2W*�/;x߹l�?�T�b3C�}~������a!i�
8l>��u��A�|�/���Ls~6q�hmV|��J)9�ì�V��d�m%Lj��p�rX��}f,t������M�d�n$%�?&���x���)1N9���7��{�m�j$w|���NL��j�ac�\n/�ہ�HBS�<-wE�F�ͤ���+����;�����]��Y �P/&�$�=���j��{�Z~�}}Y�k�+Y[
j׳�q���^x���@+��b�3�s.��c� 1�6}�d���B��ȿ�D́���pw�fM\H�?��}�!�ݓ�=��ӱ�<u�I� �������װ���^䬗��/7P蹦vF�q2������q�P�F��?�f��U�G�8�~\��W����D�ٻ}%����\7v�I���5��c3��h_�1�Zѷo.�.8O�ȵ �Sk��^|J���F�ӳ�R���Z���şo8��τ�4�V����_wF�ٽ���s=T*(j�_����.�D�ƹ���׷�V� o0��@�ņW�	�V亣�*����q��#� �c�8!P�6�+41�i��-�J	 �}%<�b���q��i>J�����������-|�\IwۄG�ݨd)A%�R��A5���h�3n2�*r:e��JcgtM1Ya��_uy��Pѥ� 5N�n�&rJ9�}�����A�����1W����3��S���~��&��8i	sນ](��Su���c�gV��>@����t?4��f���fO�Bg�O����`���!Pb_|�j��$+�
E�O���@��'�q���bb��������+!�s��֒�fz�?���XT���ȡ���\�Fo�H��!J#Z�Xq���]�������-�(�嗊O[�u[t|��v�$X1�OA���(��0C���r9�1��u�
�����&"�����:�"pp�l�s�Y!�����hZ�
�ADh��A��t8� H &���?�&d�R�%��c�3��C��FD�z3�^��!���n�p��$iXth�Gb�U�`��S�G�T^�������䌣59N �!���.N)s��d��7�ޯ8�7��J{��
�*~Ҭ9$ܐ�q;(;�^o���LI+X(�|��^%���}�����aQ��Y/���K�5���(��z���_-;��,OMɯ�'�,W���W��϶ZM2��@��&��U_/��1:Y���"Gtu��{w��J�����;ɦ��4����p��G�t��Y�Y�C���;�4�B�ˢ�A�:�T�O����5���I���T�S��ri��Ks�pg���甚#[:��,�xz����^�F�o�����d�)͠�nwr��:;�]S,Q�r)�=B�R�� �;h�na���\�`~�>�Tr���rỼ�����a�HY^�G��|s}�"���f�F�'�p����w�T[wAкn���q4V�(�z��Vᣂ�zc�se_�ҽ�`?�aey��b��'���
`Yy�����(�r��,�"}ù9ˌ�PjW����%r}��ϴ����w�'������&�œoN@�����q���U9��gC	E�@U�|衿i'EQ_͚ �����C
���~nb�u��_��.�P`s4���JO>hE��עbB����\3̅av�C�����/B��<�f�C���˳G���v)��HS��CM����w<Rj���Kp�:V3	n�����m~��(Zt��j������۝(�/�+�0ت+��Z��* 3��m���q�:~�G��~�<k�{%��샜�y��\�94���#�qP4�^�����r����#�$:�:��J P�b�;�aW��%24��k��,�B������4ׁ��q\=���.�5>�]�H��;����s�÷p�J�+s�#G��P�p��ۘ�2�TmI���(�;�8x���q�2�,��àQ�Y
~�� �9.郗�� �2�}�y+O!���h�\A��m]�@܉�>Vq�1=���FdoC5�S�����PG!D�)����CF0�O׋T\�E˝���eiqI�>� DF��%��a�|d��yw�B?�l {�NI�a��k�7�$t+u+ΛG��WA{d{x7�R������k`{"]�b��i-��J�q���N�z��d��� Grkl��O-�{�T�y�gv�^�"��I���$/4;��H@��2!���G������·"��M�iD%D}�G]�h��]_7�(|Ÿ�4d�����+w^]�C�ՕGy�?�&bAo��`ڄ���O����07溋Y?Ǝ' Z��ؽ{=�O�/)����oѮ���a�F ���{�.�r7l{�c��l���/%==(��쬢�9_�� �ǫx�4��z����7!$�tYø����;�h�b�  ڊ�j�6	Ub�$e~<�)ح�|�8 ��`�Ϳ�6�7)���8`t��X�m�We��)Pjఆ`�),m �
��+����\�,�cN��0 \z��*~�P�]�5���k.�_��%�Ɂ ��B��Ŵqjٷ���>Q������Y�_�o牥 Ms����4��<��#2y�Rm�ŕLL(��ֱ��Z��>.���pP5W�vs ���3�0��G��>��zS��[E������n��2��4
$y��Y�4��Ҝ;������� eȃ�<
bDJ> ���&W����k�/ŗ����P�;;���N�o�3��v��~.� L��H��e������=b�t����"���p~�Z0��K��wV\Q���b�e���g9BJ�Q �����i�{r���x:����z����h�--���H�C4��'��9`s��	��&��F�ǅ�ͅ�=�4HN �ǟӈg�� &J(S���.����s�����o�� �Q����@h�U_��z�����b�qK]��Y�RQ�J�Y�ȇ"�z����a��@$�Q�I�{�HVe�����@<!ͥ��+�<�j�d���T�(`|��lP�>���|�Y�3��gFX�5��jq��=�Uc�C���<�\K=o�͡����T�DRd�jw�0ُJ��!`f�PeՓ����%�s���*�_9��[%YD�s�C%����^�K�Q�>oEh���aq �n̺��k¾�3n��KSs|1�GJ �h��
U)FR͛�'؅y��M��g��Ҋ���][������֗�IvХ:��4U��t��>tq	Ӕ	\I�&�-|7��
�a��� ��H?�F?12Ues�f���HO�����L�a�}8�N�&�=���R���L�#����k�?�Gˆ��aw0��)�n%�������(�ط߸��>�V��R�}�b7{��8��ve�.2C�W���#�<�����)��=��/�I�P�S������x'�K�;IB�E�MFȽ�ᵸh$�MAZP؄�Ƚ�)���/8ƽ�uձKn:GV�S�3���d7�y�l"��Xŭ����)T�Ґ	\��~���?���a�K`��ܟ�D	}��~�yǌ]���(l~F7:V*YM�;��\�^�o��Hʹ�z�����o��t�<�<�>q��]@�0hh����*��$l
�#��_VC��@�~O s��.���pU�e��'2�2ry�������<~�H��;�GU-1���$a�3H�$�|�����j�~O���ZF/˓�WK�썗=�F����^u�X.�(��9ş�ũ�a��vgFm|���"��m۞\��@��o��CF�d[C�?!��q�X�y���������\y	_���dUu�Uz/��1Ow�B���/��!��pqa��v��It�Ȉ�W0bi8h�)]���N>��k���H���pt:��{��X6Emvx�֡W���9{q���%�՘�H��V�|�T�)*�7�b� ��ے�����r����Ũ�(7�j���?UYt�w����?Dd������!���!-�tZ߈��`GV\�k$�����	R�
,�sk� ������ֱ�]?fyb��b��1vvy�̘2�óQ	�|*��m�"�^�������x�?p)p���җ���5c�c>��J��bU�%ړ5,e�ՠ�@��e6s��=�Ҟ&/��]����_���L�d�`��,�>�.��2o_`]v`�u�|ϴ{@�n��`�h	�G��@�" �\p&�y�� j�FN �Ε�e��8w�_���CȾ��Yrt�m��.4A\��w�6�n�``������Ni�dc�\S�������H�-���KO! �X�0���9��g|��O�8��i��}�BF�_c7�F�쨌�(�;e�WpC�a,y�QRO�;	��	�8�5��& ��;��S�9%I����>�W���t.�+3}�Gf�\d��TޗT��+���\\s.���G[j�a�ማ��+6��:����k���>]A�����y��Cp�ڌ8���X�Yb��.d��=Ke�H<�� +�2��*.�>1R�U�k�G�)��c����g	��Q/4��i�	�Ԯ*������4(90\�傚���0��I���*qՆ��u��g�-��ڀ-@=�����i��؟�@Ɉ��/�R�iw�t��q�B��ze`ڜ^��\�3Ge,/F����rz�F#��u�-b�(� w����kX�
��>-�ʍ���{���%��*'��ܐ�q�ʤ"�����P���R�Z%�)U��e��۰��d��~��.׏���K��q
�me%��Z@�MԎRf�_8J��Ѽ[�$���,,�}������ |����Fiʉ3����(2X>���@@�,�A��K��P��1sǷ�Re�w���W�!P[����W�L8Y� o�4��u}+�=a��e[NN�0lݟ���a�_sܧ�!����U�iL%��X)J���y��L����y�	
���u=ؔ�vP��+�=��*��Sp�9�><���>��])���1�,8!�F���o�O1 i�v���������Vۀ�:J򴋋�/Dީ_p���9�;\y�w��K�6�7��Ǵc��)�:�)��>�Y)M�t������kk�{'�E��<w�����EqnN]���p�$q&��u��ub��}��_��D)�T�C�RΔ���xY�\"	���I�B�-��� W�>Tm�T
��Dl��4?G�&���|���Q?t�Ya�uqJ�z{�¾�P_��Iѕ�5aa���d�D�����N�{��)���"�7+��H���y؝�'�I��ti�(wqR+��.�`}����K3��X��e'xC+5��4����	�&�|	QB����6\����Xd�v,��V���vJ{ }T� ��Mģ��F�=��й塦�s��N�')HQk��ַ��x�v4r�Հ�&w� L�U@�t��,Z 1�'MBr��fFL_
�~rmd�p"�n�'.A��ՙ�}|��>�������j+��d-9Nz�����F�	e���|RNZ�S����<M#�ϰ��rA?l�^`����^�8��'�I�4v,�Φ�[r��ZI5�1��N�l�T�v
0a;�g�P\� vT��[o�&.���#�m��(+�����|���l���-��=��i��V}	_s�)1����E����
~t�ڄ���K8��Q�]�VDM�1�.;)3e��Ί�Amt0#�zt����j�����K��a�� |:����ͩeu�*�i�h��������eڜ�I��܌m;?�"R`d�������e�4i�,���JG �����]���F�?�ݧb����e��h���o22��"�J����H��_�Bg�[Vfׇ��`B!�-TR��w���AQ��?(�k�H3�Y��j 5�LpeY^Vpc	�O,�Ӻ���1R|�D��#4k��=̞s��:����L��i����6���%
,b�z�����"w�M�!4=�a���"�EKj��>��r��L��>9k�"!�H����+pA��d�C�$	���:�o�Hu_U��$N:c��#�(�ex�`�~�O�/i�Ll��%3�p�s �l�@�2���̺�}I�\���<�E��y*�W�1Z��$�ؽ��rmݩ��;L��glE�Q�6���.v������´��ê=��=�YG��� )2���>�h�e9���Z\���ig�v���<���q���7S������]���{	y��%��3�
�Pt6��c!��4���E@ga��1X	�J���RG��b	�� ��+M$c�d���{t��p�[�k\������{�TPt���V�q������#�G)߷P�:�
3�����Æv�|�s�����y����H��*��9�G-{���XՀM܅4��kr���2)���0�k�I�U�q�3���W4�=�4k{���w�E�p?g�(�SW�lM����A�������75�&��)g�G<����y�_���BY�9���e�v4���-�#�mp�v����ݾ��l�������ڎ�p�{*t�`l\0{
�r��Uh��,om)�>���P �����]i�P����`;�p};������3�pH�%-��:�!�K3���E+튏�ε띂hi,g���v��"é������^	[Y�킆���^Qc���f�i7��(�E��A�@y�I�t��4�A��;'�
���o� �|n� O\��N�O2�u�
�4�
GK��MV�K C��!Ü:��
�p��?鯒�ce%��������i����a�.m�eɏ��& E޼L0ף��o}O%�ތ��o	lt(F���I12��TR��I�+��rs�E�S=�xy
P�J��cOY�꫻�o}9��	�������_>�!��;E��m�M����o� C�t���o��S�-�d?سQ7��}�cX_�BW�ܨ"�����S��+�\���JL�����r�=��Ƨʤ@فC�p�x�'!���v-v�����|{�.�2Q[�Ϥy]���*�V��{׳�L�<$�DM=�*�����,Ӷ7�{o��$aY�����c6�
�b�3 o���'�vfL�P�Ɂ.�j �$U>��O�[�h����y�ڣ�d�qQ  nU�+����0��wJ젅jHd��YA���~�~�e@K&�9�f�����.{v�w6�\"�.W�**3(�SE��9���n

��-�H�&}
Tk��^�s�A&�I�U&��#��X�8�@�9?B6zN�N'�՜�OW�a%W!��C�\�/w�={�q�י��7EGr>��"��[�j������^��i�>��ϫ�������g��g��|�����RV�>��m]�b5x����:8J5���e#��O�J�Jy�f�l< Ô��j��������[ә�W�n�k�0�n��+kHw�Ԓ�dL֋QN_#�T�����Kc�i��q�n�oigǎ�d�p�3�KJ���!��3$:��W���ic'f���p�E�獏v����P㮀:-�p}�i��u�u��&6��4�\g �DE�o�=˫e�D%��l�_+Gpp-���~	Z}�n���O$\���O��۬Ά:��3R��|.��aB��s,f��� �`a8�û����M+��$�]UE��J�ˡ�����Uo(��K�~� �$&���(��fV�RE�gŏR��71ث�T�6����7*$�u�8B����+A�p��3��;͏��*�[�o�{u�0�k�i��Ǣ8D{�����@J����� �zs�� �\��s(y����o�zh�,b8�o��.�����b�����]!cOe�0��H��mcpO/���
菚�U��
��6){*�"9qπ���� +�|��c�Qf�
���RkZ���#eM�9@R8��ڏ:�[�����TMy�6yG��I���Մ-#��ƌ�g^���&�t�U�r�XHÙ�n�v�7��+�g�x	�E1�97�������,��u��J(��L3x��D �}����O��J2b���P� x�p����YZ�f)��vI	N�O�p�[�2��ݮtSN��[������l!m�Ս�$|׷<�wu��!n4Φ~�e"w�s�w�p��HO"��'u���5)L�6�$b�߰WJ�y�af+��7�CA�X�G�sc��r�X�eG8�������4����'[Pa��`.o�6
�>U�z0m���)}����S3p���+"����.����{�;�&��f-��{�����|�^֎�>����,+Z��}%ˌ�M��.��a��d���ex���m)���З�<Ɨa!�VT?>w��N{���g��R7%�n��_a��	���ޘ?G���%=�|�l�F�t��WP����2Dn�@`��W=�B�q��}|�_a�eA��U�GO�*�t�C*n0W�%����[}?�D���¥������P���#�ԭ��`�ɯQ@�5T�C�hi�1�03SU�v�q�@f��`-�`�j�f~�	)f�`&�,��ar�O�Ъ��b,H�`��@$���T�W�0], ���P<��N�֤��]5�v�5Ӏ��S�������F\�N�ij�'!�����aij�s&=���Z<��ߚ��H�g�j���dP H�,�hI-�w
���Ҩ2`X�X5"�x���]��$zz�;�^@��_���ٝ(�����*�2�4�I:m� r���	�F�0J�� Ndl̓؇�����n� $���}~��W�@�gH*���I-R54h[���lL9�ـ��xa�� C��HW�8or:�7�1�Ņ�JF�0��JV���6�yZ���{�ean�z��(�w$z�fK�.�%D��˙�D�Q��^�a��?�B�_fNy�wtnۛ	a�0Qgf'�]S"ar��K�g��1���Y�/ք�w`_�^���S��x�N>4���)�^�y�1�-��鑨=����O|9Ț]TGns�&
M�9B�;O����N*$�0�O�9��C0l��m�CC��!D<"����%i�k����a�a�HP����q#��I$|r���,�BۿPJ�!:D���](W���r�%0�fY@i]ĥEX_7�� ->��:��"+�5c�q]��e]ꞿ�t�����g�V�w�;���A�PEv35�
 )S���R�"#<�n;R:���jQ�
V���y[��m�yXΦ�in�S� U�P����q���" ��0,�W-C?$k�h�ƪ��`߰{0Rh����.�D\�?��S�0aT��~��ռd`�(Z�-�?|l�.��/3��Rq�m������ȳ9y$��0=�D���4mo�r�\���}��R�yB�0͛��+�t �&s;�z�,9�,�����|�ݴ������u3�x��v�)��}�h�g��1�7dva�v��SH�x��q� ��\Ӂ���E����Z���GH�y�#}�o��OZ4�Q�Q�m܅���+L�6,�JU}���p��6�o��K��	SmI��k�\Dh�5;B���&J�dN�%�P�r�M�|���<���9�}�b2��&�0=[j�2dR��!�n	2�?'Z��b�E�*!��g��\��*��`��aq3 ��F��.�g�z�x6f�I�sN�g��?��XV��Џ}9��oàQbպfh��N,��Aa���g#�����"���]�}�8��I{B�BQy�lՇ��q7�X���'�(H^�i=���"��� <�D6���6���Y\`��~ �r��<
nS���\��;m�����/�l{c���6l�.�e�»ᖔ�̭r�� ��gv��N�ob�!���}7��Z�gM��7z�E������K��O����L;#	�~=(�k�x��<�w�^��,S Xo�Kim����w$po	��p���:����a�M-h檡�^r?���$׆
\��xW�;jw+4��L8��[~%�2Ì^,d�|.��s���Z�ٴV�Ͽ�N��n��柦(97�F��	�*Z����m�H�('D�(����)@������= '��Z���p�u{�2y�'�١��:�q�\y|��S@J�m��w4���^��I�K��ϑ8K�M���٫R�[�Q���K����o�~���YI)�V-g��I�����t
���K���e�\��̝��v7�Xϰ[1O�`������+�o�v�f�T�g��\����r��+!}�[��d��� ��|~��$�]p�s-a�~��� b�||E9��C�f/�A���?3�B����.6�h[���Y�Iĩ �n}����/az4�ݶ�)��2Ib�+泈7�cDi�8�=i5|0p���Z����N_� �ԦEq���d����lI��귁O JF4Vb@�������w�6��[��gT�-bC�ˬ\������5O�i�ck�,���-0ט5M_�4�莞.�h/�0SgYF��[��X��$��%O��N-C�{tU�i��q(gi���1v�( x��;�{+�@P9&�vo͒�7n�t�I̫��ŋ��Ģ�P���l�n�ۍZ|S|բ����v[Z�������+���{�s�m,���3!�e��Օ�S
{��ʷ����`�F �2���jH-�?�$�H"���Z���%�.+$��u�X]S1����֩��C�t)�b��X��j��K?�@�[�T0w�;��������z����.`%���ӎu�����SPG�j7&���6�������Ԓ0 Z�~F��mD���"H,,����R+��gO�ͨ�pW��ꭃh�v#���k3j�#I?�Y~���p�"VGh5����C�y*��9���bd��ސ������_��/��g��Y&���W`� ��#��I�֛Ӥ�i{bXd6C_�g�n2C�R}}o�֎�v��ؓ1]�ҍ����L>]���iK�m��i����Z�T'���IA3���y��*�A����=�؃�Jt���~2�sJ�_�W��ck�伇N�iN�d^X�#���J�,T��kv��ʄ��`�C���	<n��5�{�́.Vo��'�]��p:hR=K���:��+�[I�4*���;$n2D�Қ��xH�G�en
i�"���_|��JU�b�4"#�όz���̮ᵺ#~k־hb�lwM�ز}�W:0aB_#��+��>��"ˇף��m���?���54�f�N|�D՗���l�M�7�Ґ������Y7� k�Pϗ�Y��Sy�|��8�����)�6s�f�CoE\P�;��q���mj�y������ud�ܱv�CT3S7�(V������:�m�L���*�K�r�J:U1�@[�S&� N�:E�0��W��_ ���uh2�`U�j�f��cE��m�m�*m��K_o�sd�H�=	��]���a���8/fN���B��f��aX��	\���| ���'6<�%�M�F�&�O�sr�vD�h�i� �u����V��Ƃ�F�@t�z���y��?�FBp!V��\���yO�F;Ukf̵����#V����jO�?l�D�:29@����=�RD
�Cu��U|+�N]@���0�l�af��h��_p&o�6�'~��\�����w��JBG�4�M����=M#�6�ܝ����\BDt�9)���-գ���5a)R?>�F��U��rQ/3���E�=�1��B�o���B�7?M	�eR�߱Qd��0}t���C�J�jU�S��+ހ�6J ,�.�u���Min������x�G)�Y� �o�Q��|я�c��l 呅<�	A��,r�!�dr&ϑ���&��EFr�95��1�A�F�i-�z&��f����a|�_90���pM7oΖ�dE��%��\�s=r�:���آ�>'��;�� ��$��pd�:%��>�)��"p�g���xd��%˅`�?ɺyb_*�"��S�����%��J�_�3]��W���/i�CY_yu��:pN��<����r�2?t���.&��ۉ��6�ssX��\����]����a��UE@�����dFKa]v0����@|p����̠�5{���5���inOY�uv��w@�|��<�Fy��\����_qs�ƒ��Q������+��$������a#�ª��.)t����'+%�ԛG�W�6}�<�V�KU�h��n�{:���Pu���ހ#��6�7e��$U�.��S9'�Pͳw��R2�����\�ٖ��q$f�Y��`%����D����-+u%���}����7%�-���v�	��M�(v�@@��˔>(Z3n�1�ٌ��uy�}+ףRLI��q<1�|�Zr���	�]��� �"ayH��k|�cK5��d���'§�}��9i�Z{�}���<�s��wq�B�""���C�E��ћ��t��8o/M�^V7j�_�D8G!m��dwq��=�Q�؅�c�R��l'�ι�	tq���ߘ��A�d�������c&�a��CU���v
=�|N�5H>D�ȷ���ɇ�gp�u�p��**�.-:c�t���<bD�&3��._��zM�� 18���	o������3s���C���#obe0ԿVH�g���4�;(>���D�B�H2F�ߝ4n�ʱ�ϻ�J�?��%ꟊ�o@�-����V��r�34�K�D��r�"�]�䎥+ǵO�e�7��:�<����i���e����d\36�~T2P�Q�T�v��	�G�Aw{ΛCM>�sT�c��.7 �+���8Yi�蹝J�<���Sm���ahY���rB�Y�A�ć�_:}�$�ӋuB�Ms�|\�u'��j�+q;�5�q���S�m��	:�!wJ��NȤ�jm�*"����X�.��v��m�G3�)�5I���Xv������#2�W-��M�o��Nf��Axr�D�|�h�X���L��j�����!�ǒ�53�*�5Kx�84G��u�1�^cI��iŬ�ۭ��V����w������cH��|��@d����{�HV�A
Yg�� +�g�xu� WV4�2rs��,��RJ����29�eʂ��������Cokv�֓�IF�7��`�����kfuW[��0�Q��Pw-Rq����&���h��V�K������@*�ˢr��G�N�Էe��{YX*�����K�%?�F�v�g뾘��hvƶ���M�)x�����t�g#���I�h��W�FGXʔ��J�=:-�\7柌�$r��'o�4}���~�t�B �d
?�������v�`�<�Ǡ��i�%=DYT��������& �WW�|�,�t<O9//lS�"����qi,Q�\d�+��@(�LY��R�|n�Xc���[k]*`t\��iEO�P~��,۵D��Mo��;��s����&d����N�4� �a�~�0�f�.J��O����hҊ�t�D͔�#: �j���i/�n��ujL�v�T@�����}�)���o�0P���:�W{�ҕ��:��k�~���r��%���f�E���'B��!w���x�9T@�S�aZ= ��s�qykȸK1�oP ������}�#���r�VA�<�����!k�cQ�_�a���Tz{gq �V�%���mrt͚�(p�G�D2,�Ge�uI���}�Uv�4=蛮��q� �r�>v�oV����q���ѭ�%{�e.#H�-�a �B��o/%T��r"v}����]�al�����n �h����A������s?i=��O�FTܯ�j��L��#�'���i���q����GGg[���\��̑�'�_&�" J���o�K��	9�#f�:�L⧁�!�%�E�:o�?�(Ju�4�|�au:�R��wԄV;����'�.%����'5�zK�2xJ0[���:���KF����퍧gu񇂖���q4����Mb�#�{��/u���e��>�|���X�� �(`.���W�j����~`G�c%A��
ܿ\wU�e�U�|g\c{S#%s��$$�m��F����Su+���f��\
q��`�ڌs�R5���G��ͭ܎���[ٵ�oƾ�T���]w�}�j* �w�&nu�d�G�3��@o����r�l� �f�>]�� �
J�V3�kr�AD6��bKb	�K��[�*�0a�}�6� �[�RhUr�Ձ�Zks�m����ЇÁ}�_A�Wj$��֑�G~&�ݶ"p��ò�� ���y>�e��Q(Y�疛�UdohP�B��L�d��q]j�?9�6Q�m;�r�Bk+��N���z���y1Q�g�>�!t��=����Eѽ6l'݃Z�C�^*_:$��z�0z ��qfc���I��(k1�z���#5�>?mX���Jk�ܟ���c[z�E���s�f._�g9�&��`}Ct��H��M�w�2��\��S���r���7y�^�G싢�o�iW�j���}H��-��=EB&����0:�K�bJC�\0-�d�'���k�-�f"?��VVK�����UZ6�f�,6|Gq����EB�92�����
����	,W{�z���R%}i���R����O���s6K\��~Q���:����í�oh��P�� .�bc�xQ&��������|��ᕠ��J�����!�8
�r�s��v�]@Rە\F���@x�GJ~sI戀�P����(hx�dA��F8A������>�jG����.`UDKA`�t�a
�<����nl��������F�zS:��oy����@�3Z2�����{L�{�׮��ir��E"�(k���<0ȟ����b#�2����@�~�'p� Q����ߝ*��{��T���8�z��~?_3K�|��+dV2�]i�-�[��$_���=@)
�;f�54��7{���4`�1�nI=
 �~06UO|�.�T 5qs�;"A߆e5nW���[dW� u��e�E _�]s~��n#�IU<�"�Hm�-��%M�p_XJ�o"��l7�ǡi�<��}<%Լ\$k=�va�C}����'�l/!2��d���m'��E�\�/;�N��VE%�ɜ�*�W�~�y[����/�FQ:�yl�� �֫T������*�@oH]�o�@�'�w������K�v����v�@(��������/6,���5Z;e�]�[�
��������9��#��KC�"�R2��QU'`l��K�;�'�Ǟ�\�h/�Co��	tM�����M��Q�6c8�PX>����Z��H'T�w�Ғ���G�n����7�i�{����i,���rW��N\�o�rTr��	��r,��_�/&�[s�cj��g���#Ǚӫ�؋�9�-Q�;�,���&���wU�l,�dȻ�PEk���>��m���Y���O�K^L ���}QSA�:0�� �$��Z��h���x}j��Nх�/�Ƕ�x)dO��m�biA�6�q������(����j$6�r�+�v~�˓�p�d��#����@D��:���y9+Jk��'d&�v�L��I��Uh�L������2��>�H���$wy)9���V�h�C��u��w�f)�O�ꏻy{먮M�am�"�0���N��2l�$�\=ޖ��=�C�۰�®ܞW����h�#]đ�"��c�g'���f�))j,c���Q�6P�&|�����q+*_�%��#K%���'�(n�"��aEs����EM��e�A�z��eɻ��`=�A��	)��1}4貧@�j��#U$k��z"�jE�WǊ͒d���*�h^��F�l��=�f/�]���}FgFɈ��ȍ�)b���;4,+�����G��Gu]&�B��%�����-�ӽY}��MM%#�z����S�SE�~��+`$�����"��8ټ;�]Ys�!����=�^��rp��ů�r��!����z�KvLH�3�hEث%bwDJ�YVNٓt�PD�Wy���a�?h��35�g�T��g�¾��9�eœ���1ګ�i�}����0O;��Y�me=�}���?��;! LW�v!қ
�����B�`�:ۤԊ��t<.��T"6{ʗī��u0ŉ��B��ex$I��+T�.���#oS�.ј15@T���Lv=^�n�G8n��B�gv��aJv�vů���׹*Tg��LsS��M�4�Y�d��2_`�tD��d��>�1:H����Znr)аėw�l��+~������oq�Kg��Va��p�(h��n�Aړ�@W�J�{��2z�*�h���&U!��EJ��?t�.�h�3e���K2����|fS5yC��*v#�U ��_Yw�\�Ϟ;�oD��Ĵ_X������Z��Q�
H�3����`�pr��73��9.���>�4wS��tk�w�R�J^B�����p�kNVViK�䋏!N��f$�4
"\�5U'����@�¾�c��h��1:2˱xHי/A�9�ߓh�'s���w
�,_6�~^ ����G�t��P]<H�����s�ap4Ēk+9v�?��c��˗s��/�E�)H8��x��F�v�^�'��#G�_U:v�.��uU�R��oh\�u!idG���<3���d��T���ڬ�	;u��w�:^���eO�PV��פ��e�_5G�u,2�	\�n��V�U����~$�:Rξ�uڏ4x]��N��gtc�`�:P���{x��E
y��:�ɩ,��;�xp�9�{��ܢ\�v:#Ký�'G��S��Խ�{E��������%f<�GI[}&���%�\S�̼l��Ӫ���_c��~H42�B�gi�&�ť�l{f�����v�+�i�rڬr��e��vC2Mpp�~I/��=���,�O����v��%�2
5���3UR��� �x2$<ڐ�$/�'g_P��M�$u����N~h����$��3~��/�I�n%`�Gg�nڰ��9�>��}J*�n�o��5e�/**$9�8.�,�SQܟ>��Wg��F��7^��t���f	��_]��-�z��#NtEHY��
���Y�Ȯ����Z�887�nT�v.�o ���>���P�@��=6��HWF�V�o4���8EQ���B�>�E�4��<��cD����|%_Y��A_��-���S庥Z���N��i�Xw��xcQ�b3(/wS��.?J�[,��|ߊCB�F" {'ht*:)��++=��>mb�20�BZ7x��_
�I���l9)��_�ē���74��\�Mô��YЀJ��N�{�j-�o�7����#ѰQ�'��Ҿ�N㨋HMCEmL4�L�oT$�Y�tL�kg�%+�ۂ��|A<�j�G�\�G��#,�ߦ�W�ķA�"P\K/O%c&��!Ak����9�]"����1���I�l�],N��v��ܽ;[�jh�Jk�J9D��J��{Z��k�z�����?t��M��U-�v��C��Ӷޣ���N4Ņܙ���0�sPrb~%&�����R�i�>(K�����ǻ��q$O��q�$�Y��C�H�o���}y�_��) [P��G�=�Wq���g�����^uAy������mF����[!��|�U���	�s�5a���d0����u�"�J�Z_y�9K�J��z��M�zn����V���bޘ�N61�P���`
d��6�1Z�k������ه�1|�r�<D�%�/��J��lu/�k�_�A%4�Շ�u��?"�^�bл����0ul��VE���^�(�PJ����d���b�#����?Ј;��`�*B�z1��u����q���a��f_A��9�6J�d�ԕ"V�)���tp���sg��[Ʌ���p���JE�ܘx(��&��R"�9O%0_lsZ�t��}h9��W�s%����9�#��vf�R<iD�Im���_�l)S�yM��,����=�D�p�%9��b����Jw����,h��r��'��>���q&�+�Zf+m�1���4�hz�L�� �v��*Y�&����T(�3���]QӰt������,B,�|~���W��	<s�i����ۣ�y��`�~fI�_A��x)z��K� e$+\��eM�`wB�~�ݎ�Q��7jõ�mҕ-
���� �H��ۍb��+�cixҖ"�UĈN�U�*�pFv�<K���=��wWp�˒���Þ���W�bB��!����hK������5�����&b�i�#��c��"a����vD$���V��j�Ld�W�
�X�|�"��b=��u>)�'��Ϻ�ʍ�lZ+D�����#vA�:?����4���nL��W}��8���V��b@��}!�DD��ƨ��o�1Wʐ�Mχ��ubH���UD#���~E�A� 縿u�?���u�-JS�E�ձ]�f`@�SrNf�	T������)#Y�5��!��KvUV( N3������d����F��o�"�Z7g��lv� �`�!�!��_�BcC��fQ�BkˀX�yE�������F���c)�]K�e�������"�1��q�n�Λ(p��6.#2n���Ⱥ=X ���]a��$�E3q�A��,i���s������}<Ȃ^}�7�Wp�(�vw}BÎc��ϓ�7�jh�i����� �@���&�_��VC�" \a�7ǪB]��q�M� F�i%�Ȳ.� zuXf8�6ݕ�Uږ�27�G�	�a��X�$�;J�r�q�ٰ K���+�3�mEp�l�4o�c���=�D���e_R}�[��U5����i1$6GwOW�C)�Ï��7�l�LM1@�����/��
��%�d	D���/6��z;����/��@�������J�S�H��� %nKxt���ss�$6��jBoZn��y���������m�LNA��#,�}"D�y#K%ݥ��f��8�V�w����(���|���IN�����CV����(���܅�p�5,�0���*	�E����zZD+�L���yf*�A�>vb��<V*���4+��H�-&,�����t 6eZ:,�Yڜذt�|qo�w�*�	_���� e�~|��(�/���n9�U����$��+��u�U&���I��W%��I�WC��f��zꄮ)���Ē+��LUnIF*�=�u���Gt��)�r,�tc�V�0]�EAڠ*��&���)�[ �q�.�s���;��H����b+���u�Kwȿ����a�2D�d��F^���\��n��}�C<�Im�:���0N��p5�l��Fc1�������JQXlo[C0�KL�]�G�@z�V��bd��|(��*�7�%�=�'��*�m����?֞��:��-�䉃Sy�W"F���3]/ݹa����շ��� W�Z���
TYWz7���ǜ��/�n�P��p�I��h,XCS6�GI��j���k���>��a+������f��j?����'!Z�OF5���j������h|��L�]�:���ޒ�P�E)��ɾ�u��}tרz�*�C��l�m�R���ћ?�x�|��M
A��d�Ys�\��Si�%ZF�u�7���0��^�sP�=re�P�d�L �Q܁�$"?!x"�;AKs�fJ�~��أL�Nr��z����5b/2�Z�D��C��<4k&n��aK�%L3�@�� 謣s݈y�H�n����#eb)w=U�?�e�lq^sQ�ꣿ$3�Z�b�c��l�(Ek@��"]��2ݪtj���	P��@.i�d�$�a���l%s�]�ȼ,)���}g_9�.�OI��(�����)	T����/Y�[� �*v��l>3�=��d1;>��&7j��,��?Xm������=g���'��/��.^�D��Э���M�lӭڿd4g���J�_*�ݓ�}�����'�}�c	��)�ki�}���2�}�E�+��m����Y����Ї���F�T��T�T�H�*Ur�i�l�U@$aBnO����.g#|���/7U��VP2�F��,Ĝ
����r��#X�"��=߅1�FAᘤ�kr�|����e�}5�	4+��Bziw[D@(S�&K�? ���a2����@�3x���@�&�t�׸� �s���:ʜms�4n��@1�"+\�����@��8�p���š�s����O�t/H�]w�ID���s�7��c`����|*Ĺ.uk�⭅�aIUL�p���x]��v"'���ǐ�v��+b�O���xwtES�-|��@Ӯ��#|,�������v �F�e"�V2 ��葘���7��Sc�~@��/ǚ�&o�����x}���s��a��y0����&�A)����ᯪ+�����&S�U;�PQ�*l"�K2[�Hl�&X%G�*�Λ����9$����H*�v�ͯ��ĖՍ�M�yN�z��;� ������_�'��W�$5�߻����P�D��M���fN`����裕^?�iW��e:���c�����1�������MKJ0�
-)Z��+���J��T����s݀(Nx3)��=���?���_��Ҥ��0OJ�T���L����0Gv&fz	-K]��Q�@YnWũY/;3�h�0;@�n���w�Y�t�o].�`�``V��V�#�bG<���O�6[��aH2��x`����G��GFO&��8mm�\GS��_k2����v�-]0~�<�<-����c����%O2���s4�H��uA�Ap�0s��$_}�%���f�g)�n`�1Kmo;]Tq.�*�{t��zpT�Y�b��7؆F#�s��5L�#�A�5�����~��!_VO�gT|%7ȼ�W��כk��It��]��>����,i���-�lp���d�<>��?*%���5?�*.�2���F�ųn�X�)^c@�Tu-i�r�ż�x�۲I��|x�?��\�꟯
�������5�������W<��.�j��B@��lp0�'������t׻؛���;��Vp�,�7�����d`?����Q�ܦF�4�S�>�mV�X�? fm ���qa������$}�B!�����k�����$��Ԥ���H'4�'vm��ֺ�JNI��Z�J��].%'xZO�gi.T�T�����PS�44���H�툷���"� }ȯݝ���+�s��1�M;�]�p��`u^5�$���ǜ�I��@����8�s)붡�ɕ�,4~���tT���$V�ɕ�W�P�6@q�0��E��6��r8�j���|���!�RP�������w9�����@��%,�l&�'c%q��=�P�F��s�,UK�z����	^:�4yr|| J� eAG���ӹRKG�:v�T^1�9����׻~��~p;t�Q���|Y�5Р:9$�-�C���x�]�M�9r9a�3��fq\~{k��=�[��6� �`ge���}�E$��h�4e݀�~W��=.��͢v��j��}� �w�WR�Zd�rZ�&N��l"o7Nɤ���Y�����ਹS�-=��o���l\&��J��}ШH>�`)�1���8*99kw
���prW�c1��0R6��1���%�w9��L	�~`X<���a'�Y�S������y�=�TϚZ٭��X�+h��u�{U
��>�o*��G��-n_��{m�^v|��O��-���O�#�E�`����WƑbv�N�Gc�f�7e�4ԄG�����dʹ���r��=N�����Uu<g��&S��}�k�RS𝻿�A�a]��-��b^�*;�αZ]_��.Y.�B:!^�6�+6� pI�����V8�M���)
jZh�g��d�^(g�n5�Z��S���S��dP�fN!�1��>Nl�������;���C]=�EB��fI����_FTk�{���I�X���=��ɓ�}(�	�3�O ���d�񐯒<Dۣ�*��|꿮j.��%��cd�U�tp�U�	F���+!�H�d�$��Ì�{I0	��|��]�8�k���=?&˜U�7�t��B��>>/�N�IMQ%�*A�.�5�K�"d��>���Q��eO+�;��`�T�Z���K�=̙%�����;e���I<u!�X�0c�H)��S��8�Ϙ9լU��ڜ}��aJ"�m>p]�Y��̹C�)��ܣ�ա����"N~��i<��P�	J=�ޟ۠5<��م��i��@�+~Q��C ��+k��L��j��`_4���ކ�o����s���2�B��
j�@{�M�;�	Y�F���>?�_��ecO2)��f������~��(1T���fLf����@��>��H��%' x;_kN���R���7�P��R����dO��{��QQ��|��L9�%��#�hg��iD�8���$A"4�(Ť\z�,i%�Ru���Ffv>�4A�oDm�L�s��u>����Y��XpZ���K:�G�mt��z9�*Yx�sQ�m����h�y���W۵�3[+ǘ��X���8 y�R;pN��/)#���9^nyp��!�T��,��6���G�t:OܰI���P��x@E�$�R����{b���$NH�/־�Sc+ u�*�xp�B�v[4&��H�(c6kD��r���r�Ԧ��q��R�`
xBl���M����5��|!���=�͐�K":�uPD���`���\����~/$EƇ˶�6���Wu���ρy�c�:�]���"kT�S����߫�Q��k�Ǳx�LA��7���'�Q+g�B[��SO�֒r�F�]�p���t�k'�MmV%s݀@ �B6�m�ސl��GKb�֝ο��7�%�su�*��Q����g�J�������I�L�,JP�̐'9�v�}-�L�!���-�0�Ô��ęa&��ϰ�7�.*�x�m �g͙0c�B�� "���*�ƨ������٢����60ϼ�����"z��Ϩ�!�6�/W�B I��[Oi����j#�C"�7�{�t� �9Y���V��#"� U�o޿���5O[�K�=E�6��/�M�����-��0�q�i!�� �%���&����#y�?�1��vH+��~3޺�,\�D_��40gIB	��(��>�}�����C�*z��;�ט���r"�tJTF����Q�	3Z�d���T�3�v���Q;4 �d�2�d�[�kI����x���8g,�.�����*�(?�q��nP����.��^�.Bp�ѹ��;|��e������E|�ێ����NT�#����\JSj�b�^ڔ_�0s('5�����9$~�0�3r�P/Sx"�Q&hK?���р�Z�d��O��lut,<�DB�Ɏ������(O8p�}Q�e�mg�.Ks�yW׹Y����5x5�e�k� i6cʾ��'��Ķ�ߤ�Hg�ɲp��m�f�+*�����s�lc�'�^α
���'�,�C�Z����b�R_���E����<�h�q ��k�cx0�����[-*]�]]����Zn����*UUZL�^�,�����R���l��Q���di��6�5�s���Tr$�k���P�8���!�5U�6e�H��E\f��|�� �^�b��A^a�~��]�"���B�Q����K�J���B�{�ț� ���^,w���wW����	�_���72�	��%�}fk��t8�ۇLr�ݮ�>���u���[u�Wj���hv#�h�n,kU��x������x�"���/l y_Ҭl��_������b� 9T���靐7�3
��<�>ˇ�/��0k�o�YM�3W�9ajI,:������)V�p��W�E���Y�U�?t��h�J�X�}]�=b��jF��P��A�Py1��Ii�'�&�L_�2����"X�7�C0��LL��u�	'e��b��_�܌���.��;�����;�tߠA�������|�Ea*�����������z���x����@���V뜀��/-̈́~k�����a��&�S@M���_�O �L�m�c=Z<x�6��m�&p-iO0���X]�9��O&����M��~�@���[���5��x��v����m{�E="Ou��LI&
I�&ӫM�c#�N>�;rP=��Ut��Ś��������WV�V昢s��ڕ0Xk:EG��R
�������Xz���aڿ,! �	_@,���%�\8r�J��g����������ܝ��0�m+�؞�c<��̦
.C_�)��V��OWu�:W�i��_��_�O1�תTS�j�
�A��xI�0��!���'y.݅-R�
�J����t.���b�mp��b�����!���j���j׬�*C�Jl���_���Ի�p��Z, �ᡄ�\(r��B���&՜���K8Ͻ-wJ|�Yv�����pB+n��=���}������O �ܓ��C��5�U�h�1˼���`%zL�J����2by�庈��u<nmM����웏���	��|q�#�$��Q� c�J�H������� v���� Y��L�����@������e�N��ǍoC�w�%�TZ��A��F٥�2���:+�:��uk��޷Ӵ{\�DD*�}��L����ӈ|)>�}qK>2�lշ0 q��O�����p����"?XH�~��m��X{�˪�t˫*�x2ت��u�hD\E%g�xgJfX,�#�DY6A�v�W����r��E�_�)l��1b��P����>Q6���H[�RH��X͡�[��ꤱ5�|�Ks
��B��n�^��7&m_Q|���ٱg�;06�:0'����g恕:��V�Ա�7��Jzc�S_���0d�g�0t�&_��$P����B�",F�Z�OLxM�#:&�6�U��AdO_h�Z�Sf����긻�����V��J1,o�`�5 ϙ�Ym�
jϊ.�N�!�Fh��`���z��d�i( [A�G���QF6 �ⶳ�cK9v��6�}t�?�Sz��]�ɨY�s�s��/66yz����	˔N�m����>8P���ۀ�H0���$�(5�=!�0F4+mY��ΝPnA��L���א2t?7x)9��+z��e�bRK H(��;m�ФT�@v�\�`�>r(ѷweF��WײW��o��Pf��k�*���I����0]N��{zUnQՓ�֭��R`~,)�f�6:��[�S=ZFg�mo�F�"�� t	�n��|�N���ɂ��l�I�r�jX[�KV����`N<���Ld���zwT�nht�~��s�o�0�X����sx�Ѕ^�d,:�
1�?��ຓ���΁E������:
eR�a�ˤ���W>�8�dn�w�Z�&T75G	]��������lr=I1�}+���܋Ϥ���� N1��.����_c8E��q���l1��y(ֹ��*h'/>�y��s�$��h9Ĳ���Y(�Ԧ#q�;��S�/֚il�sޥ���^+���\0i�#K�wM���7sY#��V�����Nߋ�ְ3�c��L}Y\.r�$�n���t��a�9l6�9  �K�l���GvC�"���o����fRX-�2d��d}�l�1h��d��ޡL�K�Kt�9�?M�MD���oFĺ�s����8����u��>K*������x��F��auW5�y�]o��p��!�dw�<���ܠ��d���m��&�~�B��.�Ef��h�!M*L7�/#<~+��b�/$�۽�,п�%��+9Ns�pl�j��^� �����{��ъ~�? f��,*�HQ!c�� <?=�3���bY��4���yqI��S��ۍM�{�gL^-�į�j^j���A�PUH�2q�M�; ���,)D�,ޗOF�T���{S���ĚZ���y�&�a� Q�)B�j��|�v0z4�ܒ%��M���2�Yp��R��@�ڣc���������2��c� Ȝ^F����%� 6k������*3�Q���0�M38P<��"����C
��o�_ ��Y����(�At� ˙��E�����֌|�{������@o�9���g�i�+�}�����N�xrJPĠK �rw0J��ɍ���/ҏQ`��v��+�(�L_E� ��t#��Z��s�f�ixyPOJ��D���RWa�y+]�2��ŧsǭ��s�Ϊ,3:Wp����#դ+=6��T���+���D������ϡ�j Ys���a ���,Ѩ�*�kl��m�R�
B�L�6�J�8 #a��3���#�y.��#�[5ɰ�:��2~�3��ub oO�&u�oZ3.~Q��Zv�g+��&ˌh+3Q�w���F㠡�1��M)��~r�_8���XV�<�EW���i�� sd�H)l
����BQ�dv��錽��1��?�UO��f���k�R��ۊ��$Q���U[��L�:��Q
 c�<K��~�h��i	���څ�.�d��;�:��R�}�EB ��VUh���Q�Յ��s����n�$��lg#�阨�K��\��5ݴ��t+�:dU?Ĝ\$�tɁ%�*�B_M���>c~e�4�}w�#P>W}x�nU"a�x��H��#��z�}t��C����68�R"1����j#t�?;���Îa�����I*�"�ϊ�g�&ND�l��:;",	]�7*z�ūffeg:8����'Ҡ�6BK�e�8s߻V^�\^g��n��6�ˌ�����^�ӳ�a�.�e#y��ɽwj�%0O�%iV�c?7�7
�)+�c��K������E�����X�:$�[|��^6�j灪#�CciB�ՠ��N�9B�'^�d6���풁�%6��g*�5�Ji�dB��`���k?S^f�Ue/ݔ�|�ę��@Bq�q�[��y8�hkj%��ٝ�H����~��r���.�e���D����Vl�6��c�{�:�<�( �� �ZZ�'�CX7(꤀GDnF؁�'jo��\�-T�x�6E;)��?0`9��Q1?�G�L�5��H[{xo�w]��l��^��6z����a�^��w۱��Бr�M2���.
 ��<;N � ��� �|�^������
��V����TR�1_�tD5T�T�0Q��&��z@�����n%��3e^�q*�h6�]�y�z
���r���a]���qޜ�o"> ]≚�����W'Rp��	~�V�S��� 2���a�I�LAb=�$��-��uu�0f��0&O���i������?j{�^�+�_�9���ߧw�����Y��z�[{dn��Jl�ݥ0����n��*Ϲ	>(4g�|㦷�]�K���\6<.�����z �V]��Txcz��e-nA?�G���
��:�q&�y��*�B�xq��}r R+��D�e����Ǔ����S��U�����.܈���(�r(�
� a�G>Z�{�,1���G`x=T|,l�B`���O��Z�����(�	2�"��[�����:�j�ٌ�d���L8��Z�#	�oT3������}8����i�K�2�>�l�,��z]�u�\���Q�C���x�)������x|ϕ��չ�~��֓!'N?6��*�-�z�?��~O'�����9��~hI�$�k�BjY�P\��,팀��F�&*�H��'�<��N��!�����i.%J$�B��~�=�L�>�%�g�2�<N�*����5E�C&�e¤��F1����ݛ=���$��;��$�~��GࣟkL}�M�t0���O:q[�x���2�A��M��`�;�-Uoq嚾BZ���z�=�������@ܸ9���"1�N�F�'�)���xT:�x �97��#�yPN`�bb�J0\b��^�)N����H�g-�e���2s�͠I�\��S>�N\�a>s͏��m%%�3��ϹgF�o��nB.��D3���ȎM@�J����hV�x8�X'�)_�MٕD��e5.(W
,�z���tj�UU�ۘ�:V�8idǹ�q�n�^D=�c��*�Rߠ�����A2��N�ccl�d�o���������[z�̡���{��P=��L���C�W]Y �ͯ!���&�ܗ���a<�9sل#�0�:`v;xK���ѽ�c����&A5��(��øݧD
掂I�n��0�%X�EP�5�1�&�c�*��n_Q�CY��z����V����@Bgqx>�a�8q���-�C�W���f�:*�t�í`��9��"�qr���ax�<��/�������3�+�<S�@�9��Q�������n��8_����A������7���S[�U�(W:�T�C��C4k$�I������#H��Y�j�ŷ�e���h�x�Ŏ���N��g�)����[9T���C)�y������v�)�8����_��I���]���wM�H
�n��_|����cW��H�
�n���j����>��%����CZ��B\Qc�`vv�>k����@���i��A�'y5�ȟG;Vf'm����J���u1�Z���25�3j-�� ����W<��TB�����9��t����2����3���iX%��]XD�����f/1+Z�8�Lp�W5�sE)D�a3�J ve��￟��LIC���!u��^��SJJ{�i�
��¹�2ؑ�Wv&����c j?��b�zr
�Kʹ����ɥ��D���)DHB	���ØD6uA;d�:��	?b��ix���z#;�1YR��=���^�������?Ws�*`�l��.xƕ����멥uʐ�k���Ը����{��`%�Īw���+H
��C�$�҈[�w����+����Sٖ@\�o����[d��|xjg�n��8t%���=���;[�5��RD8e3�Z�#4-�,Zf4�p���!�D�|���T��D�v��]�L0X�\˽�F$ʩP���3c�d��Ieŝ�W�c!��wG9��*'��d�,T�G���I�_�{ ��D�� DQ�����J����I��!�� ⏽D���1�Q}��~��p����۴k�\���Πq��:Z_L�-bJ�d�H^7d�i���~"7metv����h�b��}9�6�&R�����N�E�:Db�Y��c��.=�iu;�V<l�@XGi��'M�w��m{�;�>�ϥ-�J��/��mB��f��3"�����<'n�`�n�.6��/au�r/0���O{k����j3�6VA��֐�<2_�㳜]e
��S5�V�f�X�n}�Y#�Gv{�.�R/�6�f[\0ï�_��KeyP��&����?T��\+gK�9��.m�?zH��g�@�h*�M}��}���"L��=��6�u�"d��d������f�;NQ�&;�ь	���f�-�4�C�a,��,���=C>69����+X� ����E��1Bl�B�+�\~=�t�_�=��.:ț�fx����=[��`���T����c�m�4�1gïCެ�XԜw�k�'ԅ0�}�X�~ۨ�M�7뭟*x'8@`��z�pe�����*�bmK���Oy���Yi]$��f�@��n�j�EZ�|T��>vR$)��jE)�Ve��a3X�Eg�eE!|c��M���,�yH��^�܆�DO~bաȢ����ɵ�sb1��`,"�[u2���b{f� �s�O]�Ǩ�a%��Yt�eZ~��5@�qm�<�4c�>1I�����I6S������=�hę�:�U^�'-]�C�U��j��/qE+������ڎ�z;�G��a��_�ĉ��_E��T}�#�XRr�W�?צ?"w��&>JYЛS��e��Fy�b<T�����¨����84��/Sż�W�Q��/Ly+�3t���;������C��d?K3����Y?BU�Y-���U�3苻�J���ñ���v7���)H~�Ғ�No�R-6�9�� ��ڨ�;�G�wꑝ��Z�������;a�iZQ��؃Rdf�5M�i���
�N�p+�������m{J�m0*.�a�F��ݘ��f z ����~�'�*���@��_Y��F�a��Qrx.����*�JͼB�D�X��(ٞ%�-7s	ѽ;���c��'&_<`s���p6bǊ���rI�y��2W���C�yM�_p�/7)�䝤�'�<땒\� 4����D��&�@��;pE�k��lƜ��������.�ar�p;=>�A�[�+�����Q@�xx��Ѵ�E����3�d!�rY��iZ1n���n��>��lE�9�=�k3��W"�MH�|@��ެ����-m��LU���N̆�!y>e:ds�u�ǝ�$�����]���1�n��w����J�in��������� `Ƨw6���`g�7�\�'��8j��"yζV��q��َ�D0�C���&{��\"uRZ�n. Y�]I��9�S�^���>�ԯ�к���^�f��,���O���zh�@2[�I �p�h�ӹ����YǍ��g9�n��]�{̟@����6/4�/B��6���
9ɸ�R-�H����ڭ`�1�tv�m`V�U�LÈ`�h&�]}�nV&�5�Ԛ�6J����O��>8/�=_R[t�#�����N��-l���_����p�΀WǢ*Z&�-=e�N7�-9�RU~$�0�|ȿ���U�*z2I6�2�f����P�7��{uB0�A[ݔ�-˙hT\Mٰt�h�����|�QL�W!����d�G�)�-R�Ϧ6��(v���}V� ʱN�D�% �6+���-Zk5V��z�Ʃ�8j�/�Kﳙ�d!���;�Yr;1@d�m�����k��~�{U�y���5*�]7J�^���s�_jU \:��P�2����0XT�+��"s��񚑒� �D���O=k�T�gZ�{��1��ף+�_E�~�@=N����8�2��1��i�KJ�1.�ڠ+��+���)م�$ IF�s�q~B���L�M��1�P����4ǅO4�z�
��O��+� ������T�9�"\=� �ג n���[<�uUN�=i7�'GڣEA�az�_�2��Sy��"{Ǆy�	�w;�"��̩���[�Y��+��`'��W�r��܌*�y��K��	|M,���"�f�_h���<Q���r������;b�q�!&"h�8$Fb�PYF��
�(q/l������U��ͯ������.���̬H+�mNdE�#�(�3�xj:+���S��D���xd#K&Y���TF]M�f p�HKv6�����9�ތmb2ӽk<�b0�/��]�hv"�58;��;���9���|�s�����S��u��D��R��i��ׇ� T���Q��\YU]SY6��HM��ZOG�2���ų�o���]���Sq�*-rx�8�I�²��3�a'�R���"n�֐�I�L�s	S�&7k�����*^�%Mћ�d?(����t�yӕ7��w8�Q@�;S|Yua@q�)����VT�N!�:�z��<[�;`:I>����:��Pp.㾦�%ޔ��bڟ�vN��͝wI��!�~�9mI9H�����?g�p}��N)JB�mZ�X])�aȾ�nٞca7��c���[�'?��A�, �
b7�#��TĆ�~8��BZNa+���oJ^�bY���=�{*���R��xq�9�??�ϼ�K���Hw]��	 �d�l��r��A�aq��3i�! L*\Sc���Υ�1�d�[���:��Wvuq<b~��Đv�=h���Н\�g^��5n�Wׅ��#*%ۛ.���u��cz�e�Q�7X����Ş���?-���jq,�[���k��ʵ���	�<��{�@�g���cی�o��<:�냜�?�oVW8����Qh������3�=�ʒl-3F(��I�����(�D�O�@R[�t: �2��N�#��o��)��O]���5T=<:(���o�B��q��:�y���F=G��/+�m094��b��=AO�ܐL!87�K�-
��z��c����?.��^��w���O�o)VL��"E�����U�l(\�2q����K����&]����5�P�m)e(m�Dt�8��(�9%�-�X��&��CͿ���A�B]CZ�}3�I�����W����A���;y���a?wF{���{J��[WG�c<v2�*���U~ �O����*U>��3�寇��)(��Oݲ�����3���Όn���Fx�X�:��(V������.)eX���
}��T���z|��3q|��?A�wty����N?},?r;�:oo����@��>$i8��4�b{�ȋ��&�́y*u�M��/oP�E4��ZSt��sÌ�2�x� _�7�<>7!���k0U���|�3��Iۛ�[�xt*ƫྀ�Ms����>w{+���������1貗��S�d(��U�{�N�|� Q�`�<>$&��!���A��4�n�6�m��)R�ػ̱��N�v��8%L�������]�H�S��?���r�p�u���jG�y#�Aʅ��l�w>e��E����	d��ŉ|����v$֝�II��� ��<E>����'Qnm�X�R ���yq�cQ?�p�_�X�9��'mP�7�~�c4DB&7����e2K�U�A�kbW(:+-�G����fN�{0HV4Rf�I�G��ˀ�X���]���(bK�C�ɡjѤ[�HPÅֿg-�Q.4s>S_���M�+�Uz��&4�A#���ۅk�eg�je9�����o�6?��Uh�����&F��y5��8��Q��ިé�+]�����q���FK��@���]����3�J�N��� �˴d�y9�[vA���@r���(uK!ׄ= %�׆��Y���=f�j������$Koas�ׁ�)�:�> @�{M��e�W�D@��c�j�R�E�L��:6Ր�D̓7N���R��G��w��P�K�,���ZW_�6bdh��	cR_��-��)+H�(�Ȅ;� X���8J ���u�ϋ_;,b��p��윾?���c&���2��'/��/��������W�QT=~ϔd~��y�\м�[T�@=� 
�\�h��2N��h����΄#8���D���%����'��;_�%��@�e��ρT��m���c�����a�͢9�mK]�⑬�gզ�'���U]c�cN�m���L���O�4�{ݸ�5�:%�{�!S���*wN�')D�C���w��cQ�::ɛ���{*�c�����Yp�rZQə>p�#@�6)�@��>|��m�������	�eiUA&�=�,'�Fǖ�eI$�c�Q�g-}���j[T.�@�C�y�/�W|6`��`�A�?�N���
��{�xR�FV��c�4�e�&j5��9}��y8�I��D^y���]��M��ġ�8�;�X�rj����)�\�PJ�<E�tTu�a�N��I�0#�  Q������G#R]���_H�+�A�o�����"0�Z:�5��3��Z���'\�����4DÜ����m�H��&�;*��ZT�;6{-�<x��A���⍭�Pު��a3���]9���pl����rH?��$�#1���9����ֈܛh�O���!f�0nP摞R+�y u菼|~��$�����Q��~c�5�}k��`"B��wO[�q�^���I91���$	
R�LC5���*�_�Q07`#�1�sE�s@I` d}�{��2/qn۲�I��&���1����ͨ�믵�u���a`Y,&��h��^zɹ��?�Z�Oa�Ǉn,�e	����S�_ҷ���8�?��Ϻ�{�&we�m�Q�$�c�ܷ����qK�X�%�fk������Y�@c���>�l����D���!��z��5Ρ��"�UU��$�\ޏ���j"^O��<p�z%H�J�`���z�r= h���(=7986>n`�82Q����w/����z5Լ�%�Bd�k�m�u�o��r����hH�F�x�-����D���5_�±g���G����
��tYq��H��vَnV!NȰ3�=3y��_��?����
e�gNQ�Ǥ	o�#��P�ʖW`t/�Z����n�7.E�Q^����
R�����,���j"��O�-�hTPe~�k�Z��#Pb9&z�_��w����F&�eH�/�q�]I��	��nt�a�:��0�t#�j�Vk�k��oB��ߚ\����q�#���p�8��.g���$q��"�PF�������A#۽�ը�����PW 6��|N���rLsD����+�M1}�!��0���������I�8�
w��q�r���9t� ��QQVһD�Z�݃_��h��B.��ҹ�
�7܇�&��d��}䏪6Y*z����N��^S�[�A�����"�������L��ѥ�2� u�	��kW]e=j'd�tE��
a�
���(2���3犭�����Q3�(�ޮ���Vs>��V�}ֽ.�^;+z�S�J��eyF��B`��"�������Zn�;�
�����סּq�����MX@ds�`���I�	R�zY���p0t잭퉃�p"h4*�� U�,��Lĕ�
�ɮN}�=�+��TA�������\�ɴ$�^���x�ng7gh�M�#��RE�
��ە�H=�  *������AH�JkX̕��V���[�N�A��e�٘q�h�/eYT��O�Uu��� ����#�ݶʦ$��ݛO�z�3ʊ�b<k��v\�pX����t��N�YZE�6-��Q
K�(.I���U�ʂ����y����ۯ��ӄ�mJA��Y>��3Tb���D�t��|F$��ѾY����.lgZ15�Lrz���=�"O+��@I)�=����E!�(�K��&M�3B�j�~����C�
�#���$��=O���G��+� �[z����[hL2SէI���o��X�M����;>"�d���!>j�a�m���R��2٬��Նi|�ࢴ�4�wD*���ҹ�Q���U����N�s�Pސ�$�Pß("�y&����4ՁP���\5g�l�O�D������O�?	>������f��1:��Z:��־9�y���-�(M��^UÃ Z���5����ʩ'�0Y�}���21$�mcu�a?oLKlvJ�"�I*�p�Р��RR�V�-J��:��ݑV���׬�ix^7�ʬ�mOd�(�*�R�d�Ӯ)����<�0k�-<ځV�V�~��M��\q��&4\��{��?|VE����0�%���椇lNi�1B��p}�+��tğ�� ������%\m����5�~���L���v�ϵ#�zҦ�"�:�C�6^Ϙ���ڟ�_�.��HO�N���PY����ʦ#�}�>a�}�ZJpgb2,I�{�-�'7���n6��<R��fQ��4����3:AĻ�Τ��ރ������C��t�<O~�R��_���溨�oH(�F]4���W����e/�.>c�^�ܘ:�k·����yJh�u�����}�-C	S���^��J�cɋ�^������E�R3�gZ�0<�X��6R'�q�	���ZH��>��;/U�;#\�0 d��Q���YNY��z� ��-�ui`����2a2w9z����i�$�N��9���l��*�z��h�*�Al{��}r���o{��H������'S��������^�db����+�#s���gܼZ�,d<�����`�3dC��� ?]H��	I ����LQ�2+� ���������_C���s�Z�Sӿ��a˟��pEQ�N��냛L��6�����.W���K�Y��ef~M�Ѕ�1���#;R9���߯T٘�g�A c�}��	�bYƞCd,�z�/
�W�X6c[usEvY�	<;R��- �%��}�R6�jJvr��E!� O��2*�Ɠ���Q��c��йQ��4]��d5�ܱ�k���
�7u�9CI�"���3-<�w2�	�����Z�̀@���i`�:�L�97�m�qC��yu�]�Ohɨ�h�"���	D󉴐S���u����s=��su!T�s��f�9n<?ߠ��M��jD�h&7x	��7�盷�V(�.I��g{��2Jt.����ǽ�7�h%W��ׅ�o�0��_�h3��*o�8�"j����-m`?$��6���3_J=�R�Yι���B��=H���%������C�CIʢ=�nN�a�c�&/=4�� ����s=�;�V���vh�	��~o����m��0�n�M/�,�1���mO��g�
b���y�J���y���a���z/,�2�A�D���<L��ދ'��lSV��� �ߚy�kG��������Z/��	g�=�PV@������,�]�!/�M�����cU&[�}�X�-$EF�/�����o#!X��%A��T�BOM|�Y������P�qVӳ��j��*��К��ۊ�����>��^�;�~�>���\���vk!p��)n�	�e'��"38 �Z%_�n����nJa�[�u�&�u��]}��)�$�q�>��n3S����Ma��/����j4�٣�Nc�<:��jU��5����r�1L �
P����6\)�0;����k+�9ס�-X�����:�����T�8/p���$�L6�ڧ����D����t<Qi�������"?'�L_F�ⶓ�
�T_��(1'0F����e�>��)p�$�y�Y-����`��P`�n�`�Z6c?P�IhI1��Qޒ�w���DsF3���w��t��hi,=Y`�֬'��ĻtC�x������P۔T��K��{W��:QB�ˢ�H�=�D����m�����TB��p�5�٨-��ѾZ�"�BH�8/�e?����� �7�4 լ;�,�� �<�z�j��>g�Erc���W`���M�gnSI�eYYw���<�\K����^K�Y�����Nj��\� Ug6ݼ2�٫����`c^/��osyFo�`p5zboҲ���hE�R�퍢{Bi��H������&�������X��L��Ke�ꂠ��<��[�$�k��E�y�� ���6����=N�U�jvc�"�0��tJŴ��,:�a�`e�NqX�T�߄�=UA,��Hj���&�D2�e�Aa��v�FCS<��x^�Y��j�R����/�Z�͇ZcY� �5�2�1���,U����~)cu�Ħ:�������TU�f�lw���ԧ��$A��h�?]�<^Fj�Yޞ$�-��,�")��'#5bj^1RuF��A�7��h*m���g��LO��5h!J���DҠ@�򭴫h�D323�qM'��������g�nn@�l/������۔؟4&-�G�#j��-�I�5��ӵ���9��Ӂ�j�P���5����a��
A��s��+���"��#�A�L�X���v�����I;����z43��w\�6X�yk�b!���i�:+"ti�|n��::�����aEWݚ���/����i��f�M��$��&=���:�?ፑm�sS ʖ��	�C�&7��}�X�[S�iՔ��Qtt���������:�_���_�T�K�F��Ft��J�?VR߲ko�?�L�=��/b�� �&�[�DHQ!����&��4ir���G�t3������	�˸~)�ԅ(�l�N<(���F�/.��X���G6l9��꺚�K1Cp���(%��GOW�2L��Y���t�]�0΀o
�p�9�)Ε���C���ul?���:�,p�����N����vZځ�'(c�I9����+n���9��մ�����}�3�(Ɔ���K��*�[vhU��}1+�kUe�3������פ�C,FMx�n��߷22PdЃ�CM��7�Ą��`��ѓE�+Y�+K��Rq�����������ǌ��V�\�2���N�0��<u=_Ei�'�fc6hN��⢋�J�ݤ�r��\���ӻ�Λ��u�Y߹|+/�$$T>s<moX�"�|L}.+hw+�#�e8�O���
�u�e�p��f�&y[F䯐0�I�������y?�9�� �ӟb\V���;}P��f�;_L]���0��v'�&�=*Ǟ��W�p`�i�\B�$=�O�M+ox�J��`�#���!�Q�W3����ס�3ӹ�Z��Sq�I��R��:�@o��,ͫ	ቃ����l���_ARK�p�QR��5�n)��R�MЄ�A����%
�W��^@@�L�sN�%g��ȳ�^��B�\�B�'ei������^�x5�t<�/�!�㥪��7�LfE큷%w4;�����H�+i�>3�	�tB���Q���|�I�)�0'+m2Օ~y)P0�>�IWm�r���+�Y�Pd�.������Y;-6x����\Q�RN;3{����f���@Qc�& �g��`X�A'�н�l���ٌ���Wf]�YK�J��U�חw���ⅼ�hu���I��3�+01��h�y����/}�f�]Zc�q��jai#
�H8۫B������:�Z�5pY�к˷�8��j�c�Ϛ��;н�5$�^�+�L�M&��׈�~K�&V
J������D;�i�3�J�7]�P53pwW[W��1�����,��G��?r��<F��n>cg��f?>��N���Z�C@�l@�cl}(Ţcb����lW�Y��j���&kDZ���Q,��~��� �fto\��׍G>.�ⴺ.Q0G���	܀��	h� gl�{��mq���g��<��'"�Y}�U�4f� �,�W�S_�����{�q�_��X��!��� ~�~v����N��)�� �W�]���Vj�skE��S��/�|�	J�E*��~E:P�@Iʙ���� �{����8�N�D���c]i`�2���GO�J�>�g7��=AG[E���j�(��qX>5n|�b��͒�d^�*`��8�<�x��,���8�{�	��5պ���%�ꆢt��<�k��G��� [ou�B>r�d �v[DA"]\{����}Ǌ��>7�M==��#Qـʳ�R��~xހ%���7�h��t+��mQ7\%XJ��a�ۉ�y�k!��dg�]S�L���7�����1�6 �h�d�[؞�E5�D�H=��RШ�!z]9}�i�OA,sϧL�D	qdF)��MKT�����ҭ���>E ҙTS��E��<0��,E���h4'����tS�"r;��X��P{�ʅ��y%���aF��������l��0���S�	ZTf��.9�������/�z^:G;l��)�_M#�e�3���,m9͔���l��jlۭ�&Hzc���5�M�����1Z�rg����[fzu�@F����Z�\}�8>�,�����$T��a_��(��b�4.�V�idV�����j;Hb9�4 �Odz��
����Ȱ�#u�v�g'��S�0w�O1��d��tSM��ulВ��v;���#QL���'u�<���I��^5�I�+���lݴ�~�n�@�����'��u��o��s����>7��C'�/7�#ғ��M��	�&Z�SCD����{{�F���C���Z��,����P"�-�s~<�iy��%�z)EUk����f<��9 iK���~�\�A�);��k̶U�ϙ��c/�_���5j7YEJ�\j"~�����Oʃ9�$��y 1�_,�)�tև
d�YG��ު�ꅹs����jV�A &�`\7�5]+:ڨ=О`x�� 	���s�PzoQ	��ƌ��Dy�y�Spam��V��vZ�rs��]���ܷD��i��k+xe�T`#@v0��|*Z��oY�DI��a�����j4�P��Dr����='�4t$d���c��	���`����km�n��5T�3\�+�,��p�]����I��yuܷa��  ֫��]q�k�7���6��4ڗ�PԙQ�M6��<�bo�桒�\�\
r��"�A;4O�ë9{'X����ɴ�z$�hIw��ˏЕ���=�F�6��S{V�2Ӵ�R!�v/i�q�G�hEP�����i%eD:q��D���?�����}��';���� N�H��c�/@A_��y湩c"@�m��3��S%#��U���Ǌ4lq�d8n�O�h���K��p�UT�|�f�~�"�$��v
��!)�B\��,Ϛ����n�a)��c���E���>b��"
z�S��i8Z��{�+8�շ��'���,� r�[oaqH��>#l.���������v��֎��N[*�����@v��0\b79��9�*6���g��ފ%�}���Q�p��˟Q�f����\>It�w����a *~��aW/���<��wW�^q�0@�%5K�Wʈ���(��PK�ǎ�
���6�Z���uVD����(J���bҵ�p��a;�2}�E�6:���=w���ę]�R����v�	�;'�SС��%K�����&��c�w�:�SC� �ҁ���up�wɀ@�4��bn~���-�>�����Fٙ;����_��Z"��T$D�	�"����D��<.���5�i,5���ŨN�6�p;�D��JAt���Lx��\��,)�'��o\�����`[dT���4�Jf��Cp�M�{Yt�0B�q���1�@�k�T���~ߕx��F��F8��	W"�9.8��3�����U'��t3�H;�$���N׶�3s@�	��H��݈��C3X��{l������ǲyp��>g��6�_EՈV�CBb��] �`m�����.�B��Q4*�P����ޗ�R�Y�p򀙰^]0����´}��>�}�~[s%5�N ?�X��@�kR�H�!\2)dI���i���HV�0�kp�lf��t'8�7�L��<���3�����=�u.�n�t���Z�k��-aw=r��}X�\rg^�~c��q�)�ڣ��8&xq�=8�Xd<�׿ݟ�k@�b�di�p�������-`� 0���)o%��f+O��Q
6d�V⒔��eu�l>��X�􌂦�G�fx(|u*��qX��E?HB��vh!{`?%_���@f����y���6!Ru7�
'�C�7��Q<��$��h;�5v�u�+�+�e�� 6m{d��#Ie����;;����=�E�X�hi����$�Lr'�J (�~�P4/�	}�C�^U�� N��V8k,@���Α!�Gz?h�5k&nK ��֕���<ܝo7.��܍�qZ�����_Zm���Ԫ�t�o��mQC�l���xnq:��
$�Ї��{��|�nZz%�i���=�q�'��ٱ����:�H�Mq���Lf:���J���Ibݬ��5�HI��{XT?�$�������J�vv�?�\�1vٖd�V[v*f"^�o���tfX�ߔ��(e�p��6�d��6ߒ�o�e��=1a�פ�S=���K��ņ�Z�5υ�`�
���
��j��K���s8��Wg�
׫7絤�(��K�ׁoW���:�i5E�+����Ŭ$���2����G������������q�)Sz��)��%Ћe�3�oR��o���/R��k��삫d�x(��ޙ��rC�q>����-��%�"2K�uq��;
���F���d�@��L�Nڞ�"wLh��5n�	bO2,Sg���2Gkc �J�Ll��Ռ�Kz�����R����W�MQ�����{B���c��`w�X�r�L��|=��Y!�ԇ��T����E�pA�Ӕ����֋4^�M2z@���1�؋��Ι�T��Y�۶B٣$�@�65��f�=�=�Wj9N���`��ڑ�(3�V�{��3O� T�o�����{Jj;e��c� \�,;�@uRP~;��@�D�����ˁ�:��J���ֻ}�� R~o�n��4��>��a��{ˍm�'c@��3L(MHY�#���6�ؒ�1��)��%�i��pL�G��.�b��q��v�H+K��;F'����݋�	�1��'���ؓ.e �9��ce��y��	&4�����u���{	T\xog����s�(����Q`�?4�(y��_��:�C&g�<E_J����ϝG��0���-���Iy�Q^�� J:��������7?�<T��F�7�ܫ*��9�ͱ�{�Ηh��.R�� "��~ g?`��j�,*$��ǝ<qi���1evџ��N+=B�s���y��E��W{#m� �������d�o̹C�݄`��'�Djkʬ2��L+M�N��m���<�C|L�&��5��4]�J����0��J�u��d�z�ي01k��H���m�t2�e�p��P	k;��SFbC-Z,*����\�v꺽��Dd�ML_��]��V_{��f��u�)^S�/���dVW�=�	�>��
�"?�_������X8�S\���G���۷�2R�Ҫ����D����Vu�1�*L�NQ���03�7��1�c^_�c.�O����D�F�R�(HϚ�bc��r�w.U'y�
���=�ZtJ"�tTK5�K;I50�g���v9Z�Yfƫp��H<�g�J�@5�1��@dMe������T>/�+�Rto��`G�S��&o5k�i\�Q#�j��*_
�&�����5}Ǡ;lʴI��l���D��S��4s�
/횦�Z�;D�E���Y1��������L�}�6�o4|�����8T�u�6�����/�l�q��Z�����PԐ!��(��G�����$���y��~T��ߋ��Ώ�_�tW`#NR.I���t��iҁ�u|�d����6���`4�f�_ɳ��ҐՉ�f�0SV�Z�R�Lr�H��j���������dH��0W�#�p�\�,�K���)�v���p\ӕ���*K?J�����ŝ¿���z�U=^��I�PFRgkhE��3XJ��S�U. =�{脹1�"�e�t<��mй�5�~uO�E�\q˯��	��41���t�o��m)��O�biA7T���̽��3�](3ˮ��{�տ@f�5��?��=Q\��y���T��l�雕�_��zy����B$�N��M/��0��y�L-�iW�.U�J�<E�A��?�ڭ�6�łU���h�.3�]�� �Й������u�J�=F�)P�S_蟈E6ZvELPL�m��|�ؠ��������bP$pK+c?G���!q�3JN���6��G5����m�X!���Nk�0-�������a�B�6���:���߯�� Dw�;�M�:ѹ���z�]�P�/J�L�,GF�h%�^�W�g���ds~i1�Zl�W=�?c
6N�.U9�$�/�/�!֋�L��r�γ�{�\�u��E���=E�\{��o��f��D ��qw|w�X�#b�0I�g������z�"�q�&<���E$D[,1���a���"�.��U}��DP�}a*qo�Ϡ�����/� 0񝞉F�i/S� ]���.Qݸ�����@�ǈ�	��o���m�x(��<���&Q
$\U�&�P^X�\�ml�20�R�<����9�o;�/�%� I0�Sͤ3B&�Ic��K^`8�l�ط��aJ���ϳB.�JB��Z��_�U�@���iv+I����v�f�������>)��	#��8��F�3�P �&U��A���}�D�~(�5gs�vس��u̶H��)?#=����)��p�g.`	�y��\�{_����o�l��AP{^j�z! ��L9E�<�w��|'!���a7� �L7ha��A���f�zw��D���^�bTHj�%2���}�M��i?�&�ؗ݁i���w�<Q);P�(=�	�!'�k��dQK�p�k`��Ɇ�ɴc�1�E����[�8��p7���:�V*�$:��2�gl��{�3��X'N��#B�"SG�[P,���O�%B�S�I��Fe�.��ctt�8�g�x����Q����S@�&Oh�Ӂ�'����]5pP\b�>�2QFV�T�}�����ٸ<[_&����Z�Ű(��J���z��J���4�:�l5}ʺ#[<>'���cɪVL'O�.�r����/�b��2ho��Ě�H�)8��eQ��-d1쥿$��h��2Gm�P��%�;��Au�5�f�:�Ӎ������3]��]�����x�\DrL����L�Y^��u|ny��WM
!1L�A��	7O����Z���T?ḯT�|�\o=+��u� QT��H��U�n��?4c&�}�]�`�%Z�>�E��9Va���Ka�f�tt�5��6�g���""�$�.}���8�k���3�w�@Ȣӥo԰�s��c
�f��� Ȫ��OX1����C�|�a��}��p�r����+une�C�}��;�����@�2k�m�����T�0&��D݋N�x��m��p����/�I@����l tvv�׸C�b�Hw��P��n<��gVjb�g`.i��`jv��ݳ_�׻_L�C�M�b��^�B*
0�ﴻLe���Od[aH��A����g�ʓ�l�!0t_���h��6L�s�Z�#� $r��=�Һ���<��6m5a<2rU�E�:��/�?�ӱ��CiƝ�.�foo�Z"�P���02��Hmw�^ZJv2X�;�v�U�6�`Ғ���e糫�ƕ:��g��C������nL�`��ض]�A������K�"��р��U"�<Qp�F[i+�2��VZR��|~m*��/��(��M�w �%���b��aR��m8x����9tV3�;Y�Kqk���Du��`�3I&��ɯ*,�`KIӿ���-�#*��V��{�0ߎk��������-+'��:�B�XW��.�{�`,D�V�hoD��V�Ϧ�_�Y���G����p�j�v����5��.�
n�|E�8�;q|�x�~� *�尯��:c]����hw@����飱�9��d�	TD�2	�o�A�3lb�$�LU���J���� �$��`����*M�"Mμ<El� ^�5GϤVkEc?�K�s|�* paj�3����PLr�d�8���q$u�յa㛤�Cp�Ȅ`�=���1ųY��ή�t�_3�︑�8!$��V|ZL{�4�3JM�̀��L��I���{1d�5#n�s�Ұ�+�!�B�)�J�Qz,�4yX���Sj[ �`r��ϯ��Z>Qb-�FT��;l��Y��8���c��ʦ�.��7UВa�9�T~�l�<�i�*ְ|�}��"^���"[�1_T[ޕw�Y��B&%CB�.�&d�o畫��dwk����":����NJa�^F�`��q+����S�,�dԎ�?}��޴G��.�]m)wH��0���R���0t��i���C���M�PmFv���I2�Kh�N�����6%��ad<-1,Yd#��_�����\1��e�c��]���z,����*�\yV��5�c�X��t��%!��)�~��./�8�C[U���Ծ�Ǣi�'`WG��k����d|I	-�+�ߜ�nt���mo�
+;`�VV!8�`E�5�bY�n����c�'����%!W�Y3�+���E�>\��F@�ׄT�Lx��y(>-F�n�c��V��6<%=͌=A������(l��R�iE-V*Q�S��.<�0Y$����#�\J���Yw{J�SS~�]&�"q9�p�D�Ohv��rJ[�Lͼ�;�I¯W'���OR�TK��㼭t�����!r�R�����嵓�8h�.�gݡd���b4�/@izl�L�hW��ͣ�#�����H����yUU�#I��<gvЋz��7������V#M��	K4$��H��
͸ќ#��|��N �&B}�f��W���-q�
f��]�bbgT9g.`=B�G�E�<�7�w�&|Ь�J�
f@�a�&2(�R����?�e�j�{TϮP�3~��݊�.�E����a�Y^��7}�Ԇ�rF3�o�U������;�K������`S��<�]���>�vЬ�J�i��H����i��V샍��m�\]?���ǳ��v\����(d�����3ׄ
�9����BDo=�vGPX�����|����'�!��3w�V��cL��Ŧt �[#�u�d�M2Uġ�F�ȬrR&�u��"D�K��n��U���%����"��`�ߌL��m� ���ԩk��Js,��YQ�kӷ�%-!����8��v�5dl�]�]�J�dn\��җ�����&�9��D��źR0��$�uE�e��!g�c4X��;%��(}�Gp�@>o�D)��X��
��6"knߞ��q8�Z8-|G� �ޮ�/S�}�kN�5C���s#��Ӊ6t"��[^mT�[���^	�;���9�`��L��ʅ�n�ITPK9vք����	�u��rD/��W�޵^�Q�D"~����}"(��={�lg���M|=�nݳ��e���3e�i��یV����S�f���k�H:�]�_9�Q�^��,�!��շj��O��1�&�D�+\�3��k\;J��@$ӿyI[	-�S�Q1@�1�w>fuڷ�o�y��U ����cWㄳ=W>N)C\(�X���&�`�:]���kI�Hv2�O�X�o��n����+�ep~5��i��B�Ɍ�ſ�T�a.Vԩ7j@�ΖQ�#��~	F.`94+T��T���9n!g^����Ip��3��df�'��2�b�-e@��\y�A�pA��8LV̵2���4鉟�HQ�mxS>8U��8�ѳ�D��'��i)��-�e�N/���}Cޕ� q���@���2-A�h�{�����F�3x(��F�o0�r�Cw���QN1v�K�2m����n�_�O�F��L�nM��m@��[��.]�����d���_M���U�#��mk"��RK;�p����B���ɥ.�Mɿ������n�?���.QA����)�T �#=8�:�,�
ˋ��	�|��6ڎga*h�>.�'��.l�fFU����=V$��/��-O��0�$���M���Y_���(���H_��0Ηs�l��� i���<�S��R���7�)E�3&(d}׼�и��������O��$�/��z�" 7��֙;��]�_j�U�bߓő�q��G�� ,�.��~XN�(���۬8�D(.��>!x���nE~������6�ۘ��5�a��S8�Yz������a�7���ߴ�Y��]���3X�<�Ai�/�ϊNz�_�:ih�TZ��@{ۧf�F�0��u̓e�T(�-_�eH���yP5�'w ��3��Q��j9�b�n�[ɘӮa�����Xȴ����0S�iF鿽�P�'h�4e�+�!�.�u�e4,6�I��:3�5^���6G_�B��*��WMU,�2dcY7U����#9p3��O�,�
#�ٱS��`ۄT�G�!��;�O���<c?i���Y���E������G�Qݱ�
*��nK�eg���v����2|�=�~i��6KC�ƾ�q�yh<9�f�����`BZ(�P��]�΢0q`
4��'!P�(7j��m�O�Ψ�rk�B��Y� ̠�azΙ�qFl�_��5�����$�t������(���Nְd���J��a	Jg����Mj��{��*���:-�9K`g���*Ei�~�k4 �u\�
ORT8�{�`��Cyw���&�bU�ةy�����������M8��3��Q��������U��m�:��+������1�^��4	.�0\�M'Y��̏O���$O����+���n�s8A�ihY*[ Eר��&��$�Јo��R�ʩx�Q�`$�?��[1a�M���?�L��ҜH��px�t�8{À�*GCۄw2�wn(D=�9�~����$�ߪ���/��p8���堬�؍������~�zs�w-�K+Wk!���t"{!��>�E�;6)��q4;�H�k���b��y�� 5�.��[�Gy�����UKN�_�KPp�q=����X�?ڱ�u��a�'I����[L֦�U
�'p�@HŠ�o�V�_�ׇ<�峗@-�E�
0�N�E\Ů��,ay�i
IQ�Я��$ b�k ��ZF-�q�HD�Ꞃ8��n^�(�&���q`j����l���n�����χB��xn�g�c��b���'r�|�(Ai�Uu���mY�մ��� �����Z!/�ñޜ�JSJJ��TR�J��?C`3=�md6�#"H�Z��ª�8��1�ބ���,2�.V=��Q�<ӵ���o-�7l &t�gqƨ�5��g�$&�ۓ�[��+^8�r��)���E6P�Bi�b�wg�˱9���*�]�9_p�ƽ�N�\�7��1x�XJr��3� �y,��5�c�Zj��������[a����"���S"R� 5��� �o�U����Q�qLnG�HT�y���p�u\�'T���z�,O�G5d��жaWg�b�[���3*�5�.<2rdq� �؋�%�ᯱU�-\�����0F��w@rM�rZƪ���&%�N�G�IP4����8��ӣ,��\�Ij�]�{ɩ��Ǳ%�O(03N�����}���C��9N�v�ǝq}�u��[�x�<iGd�H7�]�@��!kj�J��$�͠���w˿�|k���&��%����ќ<Zd�6}���a�2<JxS��A���OX�b�C�^�U����[������,I|0�6���Ԃ�G(�S�k}�eFպ�����\	����f%,--y�������w�@G�|F�j=����M��=��C��鈚�����wɝС<T�Z��.5�$y)��7Z�D�C�~^���\�}�;=ߴL�k���$"�>��@2'�B���[/����7�U���Ah�m�0�M~��ԯ�bWz� !�)����"znR��ͷ�t������@g�;ƨ�g�>���Af�^p��;�=O/�ph�@~q�G))|	��[��eŎ)�]Y֤a�&7���~�1����q5�x��s�����Z�:w�^i3$�Jíf˶�h��M�,���t�y��(~�U!�%2�8>�Ȑa���I� ����ZB���x�Ps���M�7�r�!�_��w��V��v�?on��x��Jœ�v@�N1��<1Ra����[�#+XA��x@۳����ڹ����m�,Q�>�L��Q"sY�DX���� ���M�l�����mN:���\��;�|�R
@K�S����T�]X�h��/�;���e�"�8�]��,O�s]m�K�x*'�N�ٵ/F`f~��ՒUZ�U\�e5U�ݫ�Y)��^wC�u?��Y3;&�[���	�Գ�?�:���C0�/����c�`Zl�M�^j�xYbD�z|�\B�r�y"nI��{������N�.�.�:����g��{�V�����-g��Cɛn�C�"{c�m)�Gh���jP1�9��s����{�H�T�NG��j?��{�J��əđSq�×�|�$�m�����xЎ������}��v����^b����_���Cr�ڝ��4��ik��v�<hk��n]V�A��¬�*����1�<��*eտ�T�"���M|�� S�E	�'*KI'���ի1oUP���9��'�#ݾS"���֒U��,pҊ���5�`�Y����k�"�z�-���x�:6>��lO�mI�EP�k��X�ư� ?NdeR͗��U�h�K0c��n����kg-��#��.x\`^Y�[&���3B��ef�{�ܻ�'�p�μ�{]jÏ�?%��X+l �r��R�Gf1�.��");V��\$��Z�nk(�s~�x�v�^���묏���M,B��tz�kʨ�����+��rjǫ�
�J1Xh�{e0ׄ�fB�j�o{�O��ĥۏ
����.������!������S�_sT�=�W��m7�pζ7�0���̭U-pA2�[n����\��}��zh�����VV����dxm&��9�:�fD!誋�! �aڙ^�����T�Ԥ�n1>�&�[�1��E�iP:@-�7!N�������rt��?	��
F�'�ͧ�\����o{ub DXKI���U��P��ޔ�B��ik�P�P��2r���j�}G
Cr��2F��B*�#p	ԧ�����z<�^3R���-��n�w҅`�Q�3�P�P^.�HG������@�ef�WXk����l�8A���y��
�4h<�����<!h�| #��>�5uO�u�d��+��u��P�Xo���[��aX�%����g-A	���@p<��ӈ^���mhҮE ;�7��A��V;�������r�<��T�j�g�4)�YV�����OY��%�rʜ�O�a���0�Ω�[���
W):u���Q����3�`�7⍣`~=��PӰ���ֆ*)'_o��O��m]�{��w���0#IrHM�ƒ�m4�/�6���������E,�ף2���u��8.@O��~�V��Z9���4���w�ow�\&��=�� +��N�z���u���iC�'��=)X��E;��w���&�<|>]5KY< ��g%=5�s݄.`����>�����6�]���хv	�MD����j_(�m;:v��Ծ�~[3�B0Sɹ2t��N��/�6�E���������E]�9y����[D�R,4�ҫL�yOE�c8f���oΩK�NP�% /�������ARޮ@SwЙ7��rAk�]�Z9�~AĢ��'��"�[ H�%[kY�A�tҀp*i<,�*�2;p�:�."wuq�̨+l.��r����Q���2�x�5�V���l���Wv�����Hm��C��ڡW�į�\�뽋pZͯr�0��l�'��ʩI	q��h!Լ�\f���u�Gu�w�@�C8�#�9z���,v�"J�8�dfA{����i�Nf"�	����\�.���.{���������r��s�Ф��K�~�t:O�;g
F#���W ��̓�ߍ^Z	������i)�0����r�Z��Pc�����CH�C]���ZA H0�dԽ�nߏu�͛O��1����z��'�Le�ĸn������PiQ�qr����$ew<r)��m�D�Q@�b��?E*D=�,�r�E��k#/w�`��:��š�6��ɼ���-V]�ӭ��Q�\T\���[�� �M�B0H=��D;r�c��}H~L����$����ݗ�uˋU��ҧ6�j�� �;��h�����T̖T�$�M�ѩhRH�>��̜|�2�!�4����,_Z�h��9�o������eF�n��ꬤ\���W����%����-�/��C�pf��-Oݻ�1�Ai7�|�p�l��+$�s�b�c�{��4��A�L��$O�B����q��R��s�A���(x�rS��@�O�|0�G^��[k��򡟒�:'_�;�#wm������-����ĘQ3�J��'$~�_�\���J��obյ,k/V#��O��H�Q�>�U°�g��A���p0���SKZ��ޮ8V�{n�D0q�#_M�C�� S񝻲ؤ�������e�4y����{cdL@W�TW��3�p��c:T�-�����ɡUJ|#�6�zU;���`3Ȅ�T�O������`;^�s3Ԋ�bn'�J�q�46�.@*��G�#9����3a��yuԪ����E���Z�(.f�KQ���:Lag��K`�}�^+��x�&��ډ��g�o����ǔ���Y��㤀�'�}��T?h�E\�m��a�UQ[��F�|�SD7(]�&&�P�M1�3^Q�O����p�\��\�3#���詧%v١�h�	.ڂ��x���9T飷CWY���}	3%�ƀ�7���%�Q�=�n$V�G��jM�0�n{�T�]J��H6)���g�`/�N��ɛq�e��F����+�kҡU�]��bqky�C�q.Y��%~qx�|B�F���¸�{��i��9U�H&h�&�4������_��c����I��M׹M���L� �#�ر��F���=�� Lc»��/���qI18�<"�R�do����z�������5,�P6t|j��3 t�Gxs��w�}�3HAL����X��I�㢽p�QPR���u= D�2�+1�=��'�{����n��������� J��[ZΩ�M� X>��� q�lx��Q��<��ԉ�^�%�#�;��g�	{r=�F�rF�*��g� �"�a�(�pf�֕�B�'��g�H(��Lm���l��Y#�w�ːW��7����B.�FQV����t|��<�+�^����̧�_}�� ���5���1vզ�^�3u�y'!�u��Cx��+�����1Vh���Z�Z��f�$-R�f9[ܦ�30���;>�������x~�zR��Q�Z���-���*$M�%b�D��F��l��
�CCzw4��.�;�a��!jPD̛+�2{��>u-�y��k=��ԣzm�'D���A��{���ӅH8ߏ����@i�W���� c_d�5����3�H��G����*��өb�5��^��V[#-�ĺ�/��_P� JQ�)�����qR�8w��Um� ���q��c��>>� RC�|7(�
�@��>&7�����Va K��(E8n�����n�u�pJ쩽���8ŧ�X�q��<y�|�H�Z��+�M��eݜw�Ujw��t���aھ)�rI�* N��q|����/�'��7��ɉ2�!�r[m9�#G}9�Z���J_b�)���;���{��__�%�E�x^,ݗ1/����4���X�q��O��HL�5+��'�=��v+�m�r �+u�C�����Ԛ�9<>sv�YvZ�y���0{������]8D�=0g
+ nҘ���B/)�Z�O�w7�.�@ؗ{����~�p$�>i|� ����p�Ep�6�Cc����
�׺�~γ�Y䛲泗z=
H�'�V��F9��� \e��`�)��mX�Y.bQ�Vn���'�� ���Wi[�P�v���S
�3��ϯй�C"�����q�Xƹ���)ܺE�U�����;dH͝�Xcï6�{̪��@@J����<bo��	ǛM��%�OFOF�-��	��nj�}�� L�s�&=�|$�\?��@ٷ6g/c����2�P���
&�Q%���!�(v�q�a� �L~f��i�������4�0|7f(������0݄�=%�ԭ�-����&WlP�Ez (~O��4w���wf��F`�t~�˧�δ�I��|�!���5�?��zO�!L>�;��V9�Ă�J�}O����o��T��?��m/
��"������0�f �%�  x?��'d�
��������p��͡v.�J��p���81�D���q�r:[>�W���|;�ݵ����M`�vdi�:�k�iX�E	v�_m]���Ӷ�z���F1ܩߔ�������
w%��X�h%&z�W�yܖP�e�L�p�C��vE�av�4 '4�p������ ��X�W��0����x�ן�ψ8@�U�w�ܑ��`�	F��I�������-�o>�������Q(��I�Ję�y�8�z�9#:�.��Z4bF�,A|�o��N�{|�/��&j�ZExxV%��4T��~����#A���9��a����&g�i�����R�N��G� �gX���s�q��Dҝn�K�zg�]|�w�W�8�neu����h�'q��7�����6�� E�)�z�V��@_��=3�� -�K:YY�ͨI�cOYeι���
)�H��"
��>ɱ�����#�\\Z)��ͧ����G`$��e��$�r���
?BD�ٺ�˶<_s�	���P]f5��L��!� jFi�Z�`F�0�$K�Cޒc���>���P�t^���ryO��X�P�3<e>Э��Xl_�6`���9�v.�#�d���ӧ��0!��f�{�J��8�=&��\[��x�����*��>y�D߽��GseB�V��W9�oL~��xl,;�p�AZ� eB�@���].�g~��I��ߡ��H���Gr�B$K�
�/t�-��9։�IC�?����Ve[��R�X�y`JH��^�sF)BOa�M��
�(���z�B0MjJ��"JkԂ���.�i�E�}|^���:{c�.���'���*��DilE�mT�x|i��HU,wQ}�ⶽ�I��5�R����ΰ~v�-�dh�ZM:$���u��ɰem����g���#]�� h~剪<����;����D���4�46�hkt����M���o^���l`͕Xg~΂�dW�tX��39x��%�"���ig�K��7@%.d��a�@�?��OJmT��9�9>���i�Sj8^�̏��]�֑�F�< ����l���7��@�=�Ԇ��?wu�݌��	|H�m�*���^_��K�x,�.��c�h��L"h.��� �g��Ls�S�d��2g��>=�s�yL���#6�'\m�@!C�$�|��$�Ԫ�U>��{����I{(z�3�<��d�j����"�|D��^��k�6H��I��Y��g4if�h�!C��b�MУI\�kQO+�W)�S�w2��o���=��m[��N����������2��U态M��Y�&8���ڷ!W@�KV-A���}'���ɖ`8�䈄oFf�2�3�Z��[�8����:��>@R0���q%i9pM־+kgќ}t�{vKY�逝^Q�~q�C|VAc�{O���K4n�2b�$)k@�z<e��W2#��`6J ��4�,�����{����&��{�`h���ihޠ
<�t�ߙX�x��k�T��9�����4/��wy�u�G� I�{^Y�jY
�1���22�̠��J�u�FpA��i	��^E^EPW��>����d�؟+����?$Du��V��!=����։F�l]�So̔��𭁣�jiڊ����*�z
�t��c]@aG��S�B%2�k�:�^���;z���-�<��0��$� 6w鉼P[��Qeᨷ�"*��&Az,���K�@��~Ԟ�nyZ�
��G�臓�����>+w<m�M�xwн���*lG���x���hGfGg��42o������4�08r�'_Z�$Q�������ҟ~��!�y���ZLzU:�ؐ�g��8��W�B��]V��#K�|Q����P���Tm�@0�㭾vS
/���5!&��2��˶hjy[���q�c	����H�Ig.?]�Lgz`�:9���F��j�M�`�m%�y���;��-&�����5@�]Tf�S{���W����ֳi�,��0��%/���c�'c��>�1s��v��M7�0M�j�
�N#��z� ����O�4|9яSx%
���h�m�=r��`�5������?{^��&Eü��F"�`,9
����D3-U�.y{y�g�-O����/��Ivj��1��=���7����Z���>>����@ΰ�h�WA�G6r&7����1����u)
 �C����!�_l��	,������(����<��p��	=$h���l��D�	�g馁t(NM_��r���\��D2�.�y�t=�5wD�Y��w�x�B�o�dַ���V��$�S�joڇ4hd�_Uu�Ian)8[�X���r{;ebK�*6�y
�c�+g���3׬�&�q]\����G��6��Ǖ R�$����z��ב���R`}c���k(@��E"~�� �{��б��eo�U!H��2aY�9�>�%�.@��ja�r�A��a�k�.2�'%|\��B/�o��o�9O���!�h�~�	�;���A7L|�He#��l�י�xG��/�p&z)���ED�&a�u8���;���vM��jF��Y��{:0+ͱ�

�NƷ8�K�\�-�$q�\z�ʭ�b��?m�u1����W���y�"ǰ�"�7<֮��Du�T���-uqdj=�ܯe2�6P&H�%�?��&ew-FC�Fxx��\<��;�	�S�u]n�"��V4ֆ��>�D��d�	���n�u���'aթ��3����n_�h�<\X]M�)��>���n,����V�S�;۔��uz������ �/���X'jFw�'�{�x{GR����Q��- 0	o��u(9M	�$Q�[0�F���P��8�D��:���c�����e�c�B$[p͐Pz<����l�D���W�Ѣ4��u��R1�պp�`h+<����<���>�*�8���|�j���2��PCt�C	��鯪�^Z�5���.ά�r>��(HJ�H�-�f�ZfN�����#��x�-�9С{!�&�ڛ�>Fs�4L]r����X�Jp<���2���?�i+i��d?�������V�+���HѶy�vhP����%�:�e �����6JYaJr�b&j���:q5�t�������SJދ2�'4?=���K#��^�R�N�W5�P�R��!s�B����v�Mr��2,����gz_�������r^%PX���&Ó���о�\��[�G�`��e�Wۂګ��h�2�q���X����S��`���4&�T���נ^�� `�6�����t�|9�"�F��Jbi��%��ã��;� ��u�W;�VwSk���(�$S_Mc�ٔM9��T�/�%i�"���ksA?���OZ2߷�4⥉��$�6�eZ�T��$���U-w{vݒQ�=�V�,�[���f���^ȣ��*E�F��Џ������:���G�Q3�h�F���Sb�{7����W�[�F��2+eR@E�0�����!x�V�Ta�WJ���1��J������i�y2��?B�`,<dٽg��#�	�����h*�a��ϩ'NfA�ڙGV�&p�D|h�`����8Q(�D���1�"r���0V4����\�R�_� �h��c���n���?QV�����1k4�<�Zp��-���*�:�:����T�!�.���f��˫}�jL(�x�l'c��	�"���b�羡�l���,�/g�d��

�}&C"�a�8��g���b���ǐ�}x���#=&�i�O7ʫ)�M�,g�r��k�����'�2�0�[;��`]�}cM����E��)>���ԏ�)ݏ��Y��n*5���vɽ������H����9=��n�xv��W<}L���8Q�6��E��N�S5p"\�m.��%��8#�;�Q]:#��b��9R\[�>k&1�h�M�Ԍ&"���G�<�H��c�=^��1h�e�����m�d��Xa�&A4����:azrrAz��T���rP)/i����sq@�T��$�TY4����@�*Kj��D�B�x�"���1��ԍ��!��\A���|Զ�����.t����� n�kj[��<N���YI�"�V�%�e)k2T�E��1�4Y�t5��NL�Y����3�y���C�V��y8����R��	o"⚣�H⚦1;=��v�J�ף��Q�:�0C��OZfDA�S��U���d��uN��)��]�G���gI��
m���fqW��D,��o�SE�E)��J�bޔ���'�L:z��kE��
7S�"���$����D���3���b�&�5�;�3JAM��QJ�2�i�'5^)�ܰ�mD\���W���"^�kbк�Q�H�ՆV��t3n���.-UCs���<��кm���Y;Ӵ�����B^9�+�+�4�-Q����5������Z��a�#	��Pfi�o�[t��{h~��93H��
~z5�L�=i��*Km0a�](��,��knV���v��%���2U܀g�d»�ӑ��o����R�$�(����WdA�#��d�O0��>��k��_Qe6rW������)l� [�l��c-K��"H���8z\�bW�4*�X��q>�)rWE!��%R�>�>��	O��|��Ol�U���`�_��A��1��̄��!3I�ړ��#�<}��z��.>Ye�Q��&�lYy.�";zţ�)׻G���&�I^d.�(md�U��I�Y��~��Y��Zs�d��LJ��������6Y�wC�I��&���FM,H��s�5_2�V���!�L򡮆�5�ė�GI�F���k&W�G��K-���K\��-���o��롵os�?��f6R�H�~@�t��jix+��A�����M�%�po�����cia�x�u�r7����o s2\����L�/�>�A�zn��R�?.Nh;X09[%N�\�ew&Șh�C��`��؁ݪ&�7�́�)�0�켚(�a������5���O
� �Ɩ{�Ȓ�L�M�ή������n6��]��U;]��m���nM��Di�xC&��������l�@Y���G�p�J���B#f�j� �mQ󠡺�	r�ڠ*r&B7��K7���d��G\��j	��iӁ.�;�`O�����s�pU�E_W��j�$�,{�W|�ڋ�C�����d7<�(�ZJX�[��(�)!Gzy�>o1����<a� E�����j%�)��A�c��vZ��W��$�g�nf�
��C�w*�[��֬��@c���~4Cu����ǎ���7���i��>}d���Fo@(�Za[��Q�*jO#үt��-XZ ���1��yG����Ն�P�E��ː>�9�`�`1���㮫T��/��4����N��=���w��$��Q�����1��I�k����
������Q?��י�9��k��4�N�eԱ�����0��vG�8�S��OV���'���ՠJ�9i���v+Y�і����Cz`Z��nA��)�"ꎂf���xu�$S�ߧ��A"f��&�P38��V�O��=ZQ\W�o���y�`�˷8\	�@8���ou�W��Ć���`5��O�����Y�ش@ 12�)��ᗿL;8x+;f��u����1����'6a��ǣ�[�����|�OGU&��� ס�v�Bw;i8=��|�0���$�W��46����	]����?������D"�.��<|~\���0(A�C��<U�/J���$�ڹ�Y���1��r��u�#r>A��L[���Ɋ{)\��E~�[���=��b��	���Ix؋�'*4Qw��!� MXa"�Sv	�0Ƃ��#3`Ym,�����:�/m}�;��i��onG&L=�z��ޅ���Z�غ�A\!̩<k��./�
~�|,Ui��N�j���ōN�]?�mNe����J���f�V���xla��`�*������2'~�Y*�sP�!�2s�R :����Af[�3��_ ��9�|l�Bz���R��������#���Ux
��8�C+��w�^���X��F��+J!�<��0I��7���J@^K���p�.�]8�d��sG �O>r9�'Z�-�]�N���Q���t��|�M�־
s���lV��,���&m�$]��Ϭ_ܚ�
k�k�;�,B�_��.L-b��j�����G,���@�rf���Wٽn�k����Ӎ����Q��BX�����,r�Qhh�l���
9J:OaW����|fI*��e�,h3�l�����D� `@����o�0��Yot���*$.�Q�F�az"�<!R}�B�'?���)�ڙ� o:,�~��⤀c��
gtoF��'��l
�aaJ��^?TO��t��l���+)���B<�A�QJ�#Q$��d��Is</�u]��d/�fG�d�_��ձ8̥�b
̌�Яrϱ���HvF�Bߦ&�_�}�M�k����g=��/���Z܅��&������G��v��RI�>�<�����Cs��.�=��ho�L0_�>i�z~�nm61պ,]^f��@$EP��P3�mf����Ǯ�m�r��>ƟI��׶KKi� T�Q8��qJ�S�nnv{O���4^�5�H���Y�X\����M�sg�q!%8�yv�O/�ed�PX]iT��k��!�	G0�r��G�x�� 5��4L�"#����϶�:Q�]��;�-p>�G�6�*���Q��{�^\���d?e$@�.��~�'���mٕ8�a��"�C�-�t�!@\"��|�b��Օ��g�_�(+�|k�Є-ń��"��X��*����8��:{���Į"�C�e+D�&�"���ao��$:�����O=�#�T�JJ<���e`��>��,�����ArO}��	��~U��Q��ߥ�����E�f�
��]��-yY�,1G0�d0�L;�쪴�Mϋ��*�)�'"<��v=�t�=)��#�{���H�����Յj] �b*��H�4��8��HWRx1��`����Y�VF�5�Ĭ��u�M{�:�5k��9�I���9���
�Z[�Y.�pgrG����Wd R�P��˿?뚇+Q��B��.�%<D���Q%w4�iA�FW�S�ԏ/��p�?�����2b�������ί��Ӊ�����>�����1SBN&*��}� �'�D�B�Q����z͸t�O`��'�`Z�U�7��HIO���І؇��h�Echa7#�����E?��M<k�5^^�T=������4O�b��`�P�I4�KI��6��m���>�@�p�3T� �,L�����]�XU%T�J�F��9�N��T��ʐ_}�~�ʺ�{<����=�.I��^:���/�&��5x�D���󷾰z\�:�p�!ъq���If����.ͽ�/2�?��+�����V�������&T��'��OƠ������(AS�!���[v�7t��,k�1�v@��J�;���]E��Kxm�N|�]�� �0!��63|L��;�r���i`�'��}*�%��)MT��)bvX�)2�W����YS���:�:5.�(u8J.����|����/ј�<������i�n.�C��Z�[���r��p�r��"�o�2(���g�r�f,l��s��Pyd:W�ୟ[��yZ>��yG���#t���xd^-��#?�9	q��?�5(on���j���}�d���&v;���q�`Eo<��o��F�CB���#Q$D!D���Yܬ�ϒ�^�X��zF1�Cw���X]4g�1� @��ďu>Ж���螧�ˮ(�#�5ܙ�+�l�\�����xS�ɑ�r�U��3�'~�]��3�S-����v� �&��cj��H@F��	���������k]�G��|YP�te�'E։�ҹ��=펷���IL�m�Τ�U8<�b�{���%�4`rr�u}��#�)wu2��hɠU��������eB�wp��� �[����\p�2#/`xFs|�E|�qas�޹��o���|[���3�jKk�:�(N1�ʲRP�*�A��q��w�R�%�$�����1�U���, #��z�L�4�ܯ(fpA
��1GI��qJHxϞ=B��i����
��ܠ2�T��#ZF�������xsv���e3<�2�.�v���~�rx�Thqkk[�Ի},��1�-�b��ڮ�'�O5,����̛6R�S]���}%�Y%΄��5}8��U:Bi'�e���2�pFA���[��hi�z�m�=2�ԧ
1kL�d���o��8����^��	��O^&;�:��a��[�4��[�k	Po��t�{=��X7���n^����xqf���%�5D+�cT?y��JYgsz����C�����5�\I��ߤ2��5�"ۋ���2:󌎶:�0JN����bCl�Hc���!�iUt����>G7c���@�x�_����98eڧ�k����������kbtX�V�������9#-l�P��ድsJ�/\����c1lR��RP��-��i�	��g�M_+E��d�vtSDi4�s��y�W�GR�'�q�vu�g���l�Ѕ<nІ� ��LD^�h��I2&YxC�0���R�tC%n#ku��Zv/�8y��J�� �Zٟk.���@=�y̝��H:��yV���:��W�;3Sx�}LL��������}Cv*��RF��E4�r�r�xFJ;��ѺP_�ˬKn��-.	!�oơq:���a����I���HKb!�b�,��_�?����zd��K\J7��j�}���p�r(:/��Us�A%����83������-鬮"4
Q�q������
u�����i �w��ɸ�8��.���L�P��H#'j@�>X��{��"�w�[���B�)�M����N���޳�'��^��O ��-^�ފ2��D���m��w:�	�	 �6�����1�r�S��B��m`��";!��hE5�
w�Z��Ls�8�v֦J�=��W�D�c"#�s�P�~�ͯ��>�\o��L�'�U8�4����j\)�xyn��B3�U�I���Z4e���-�(���gS�,2jj	o[m�t��9�͹l�Ã����\�]R�z�v� ]����Ib��l�I1t���+c��䅿��Z-��DF'P3�t��sl<[�<���'���Ü�r;5M�0�e���dҪ�6�>r���h�"�kr��W��ültX&0�Ҥ+
S����B!:���S���{	Igj���pYZ�=TxU�)��W�7�MG�7��Q��%��ӽ�np)6~(#ǳd6�4�,)dm�-�,�o�a��u��pd���ܪă(����cWV��|�9l�ʧ��B�6��V�,�����h;<T��,�&w��ImU�P^I%6=r\AU(����ӫ3���$,��j$b�&�,`g��(}�bܝH�k|�e�g�5�����秊o��\�I����rHK�ߋV��(��̢�`G��Ǯ��� �mm��$����|V�����8�I�:N6���[�K5�;���_���_�3]#�"���>P�D�r�2a��͇��6��I�o�����^�c�n�J�� ��k��7Y�܋/�+]1������S!�%����{����0'�	���5׃ڂ%�Di;|b�NB݇���':#�&��
xEM��)�� ��J_���Ђsm�`��$y֝�G��$��,�c4N�	���ѐ�����&�L�N�W�PGv�Mk-����7 � S�X�3?wP�DB�z@R���Z%�I�'<�3�{�]X
F�u6W;K�ԩ��Hcس#�E����v/H�=X(�׋�M<�I�aA�vk�^��%�J��E���� w�ې�\֛�E���%oǕ�1�PQ��jϫZaԙb#dͶ�C��W���=�S")N�ҢBģ(�����R^���--��oF@���JHZLЁU�N��F� ���m�
��c��,kw�r�ݬ�Ƭ���K��x��NBnJ�l���-�E�_�}����B��`@	���aS[2��n�3 �Ǟ6q���kd��Y���0Z����&����9k�����'���w���г�^�Go]ь��a7���=�Ζ���s�D�w�^^GJ��|M��ǿ�ZS�|n(C3,4���h�:���ކ��s�Փ_�7�x��9SZQ9����3 �L<��}��C�r'M3�j���N�n᥅����f��}��|�'��Vl=��G&���2�Z
�le=E�6��������>���h_�/�HئV��(U픱s�:# �`�"ˉy��:��-'Or�B��ѐ����(ES}7���@��0^/u&���I��=X��#�W<O�C�_�����.��~y�t��'-I_!����H�_�����$����;�*�hG��D|��f��tZ[|@^�Mv�EoD��l�2(��4c����z��]�(V�D� �v�f�@�+�$l��ꌑ4�-��^ۃ1՚�<A�e:�&�;D�/��Ug?r���j����F�s�Zٴ�F���vE�J��H
����v�R65$c��c���,??)��S�
��`��E�����RJx��\d��V��#J0�Z1<.�r��h��Z!���<�i/.+��͏�eO�E a.挛�H]Mz��!�a��,dn�����|���O��^(!z�Ȋ�º��#Ew��ֲb��I�t���UK�	���h�G&�'n�>�rk1�3H��_���Kp�6��jg��cM��M��r9�����H�YF�����4/�}JIR.hN�P�����q�� QM�#��ٸX�t�7"f��k���L6�� kV��zA�)}�V-���?�pƅ�b7gZ������}���C*ʓ����xG�q�Ɍ��o�ƣ�ٛ�\Ȱä�3F{%:�U�<���x㸢38N�,t�f �Pd](�ʎj�J�j��E�|���|sM-b;�5���2�����L	�s�G�kh��!��s��h��>d5��V�
�Y������#G� �@�(��$6.�|����Sv@�۝B��hyЁ.
��'(uU�M��i�M=�\}%�(L�8h�\=������m�!�S�:R �z����[���J��ʝ E���sDE��Z(�`cS$C��ߖy$<_k�3[b?���z�n�F�x��S�]�d	%ݰ��+�P��Q�A�Bx�א5�=�9J�:��ڴ�����Ov8���$��AI�X-�h��������Gy�>��:'t�l��~�bvF��Ǖ��N���a�Ik#5 �Ɂ���I���Jӫ4�L����X���je>'�A㾈�$�Kq��}�Ob'���-9��C�gHw��XQ.�N`	.��Ǭ��?���٧��Y AC�eɹ\Ng�ѧ�	*�Qc:�6��<�Y]���S��wа�w��.��&j�=��UC��6�a<$�� ��S��-V�7�T�d�+[�<��7���q���'/�5�0�'�������V�?�h���y99�<�4��T�x��W�vB���<#�G�#j���/��-AIsGk.-!�jyT�n���L���}J6��Z$�ֆQt�Z.�	ht�o$��L*�����e�_)��t-ErvJR}�8z�C��%Da]A��;�<�����/�s_��-^�5Z{*� '�.����A}y<��e"�����n�e�aEӝz�� ��6΀�˟7���V�r���.��7��_Ⱦu�^�ʺDG�h��\�W���x7)�l�N�0��Q�Ra(x��>��K41�"�r�c�� sP0��!!���;cK���-2�;˩J���|J���Ĺ[Η���+�z ��
5��F5�ْ,D7�\����c	��X�
|�O<�i}<��e3���Y3�VS�����-y��p���?�9&�ͩ��Y��Y+@�}����#��������Q��~Ԯ�����q���-G�� ��  ���>ƺ2WHM-&�����奛��8J�#
[<ߊށ�1��+�1�}�.�k�/I U��R�u�)iK
���C��Kxg��K�������t��b�h:���z0\�諆��ad*bs��.��R���_&{y����'�
'�ί���8.���B+C���5|��v�'�����-�{3�p�����K��q[�J�#_%y,��AZ����p$��U��kX!=N(ҙ*(����t[�a����3	��&��������l����nod�i��,#�?��Vhg�QCA���b?�P����x�r�=V��K�Q��1�8�;r��~�4�$��ɝ"�F�� @��[��P���_�F���<N�p=�ȭ|k�j��-h�ks�i��z}TW[h_��5�M�͓���z����;��ڗ�po��|J�!�OA�^Ϙ��>O� =�@���wT�����8�uE`XZ�r	�����,)��e�r���!?�]�E��<�i�5A��7������=ۄ~�Z��(��/�4��I�����kF7���U����Z���\M�Sm�q�c�A�F��]�]�i	F���t��\;M��l�f'0��聰Fx���-�+.	��(��}6�Fq:�]M��q]�_��'I%�k��s�z.k0i2�әt������|nJ^)t8`)_����g��=�'=��)�ﺧ',��O"
��tv)�Z߇m�4�g>�T|�o�T�e�e}m> ��1��(��LЄ�5���{qd�+��{<1��R�)\�#� .0m� q��!�<��{a�Ŋto�4�^�cÒX@85F`�b[�
��+�'����ۇ^�t�l`�P�"�Iѐp�#��Z�߳�'�%��7����&��+����%g���GRj�B����; UZ���(_��J��H:�x��~��v�v���_��е��wb�zΓGZGe��:�^�^p1���a$QCׅ����f�����+j1pg-hө���D뢿�CI񹛞'��M^����io�Q�h�f3�3�aצE���=�\�`��r[B�u�ǋ�
c�׷P<{VO2�'�0I�����9��pX&�����ے8+\Q��\��r���,�
5 y@�M����*�4�u�""L?F>֤c�`�����A�!Y�ȐK��ӓ��c���
`�F@�.��t��d��'QQ�v�
�e�>�7���)q	�,n���t(����U*�Ύ�.�-�����6�
�/_���}5CT$���nlh`e���&��e�s�z+�ӊ*MU���+7� ʓȩ���=���f�%�����P���ņ����E�\���.��S��f�/��p����)N��!B�uՇz�#�op�M�~z�B��̋�	 �V3}^sX�a�w��QL�.63�=m������l����PHi-!6�����.E9yj��+;jF�ِB]kh;hJ?\���B+�l
i�!�����󠱺HtM*�1)/�l��s�-�{ڒ';���p�g��M�1c5�6�*!nV��>xg�f���9��umHl�-@�ʡ�Л|q�\�{@'�[a���ST.@���+�y�5�ϑ;�4�AvM��n��93����e�M�	�uV�jo�KA[��5��3|�*�C��65�������t�	�QQ	8Ww�k��Bڇ��s/�$R����kv]tt#��{�m�F!Z(�6�b]eLB�U�5��W�Y��XI���a�>y�_�w(ۈ�d����	4B�)J���������#���P�	���>��X��%O3�s������V"oÛ�̣���X&�_dv�ўd`�I���Ut d5��$̄��i�"*tИk�Q)�z���PZ{��G�/����!�4��W�<��<�5��i��D	;��qD��ck9���U�l�0	?���"04���1���z���4���bҕ��Ӗ�7�.u�������`g���W^��OUp8��BF��gS	����f�&Ԍ���Z
?�%�#��+�($$ͩ)��B";��Q3m*��d2$�4�=oz�4�_���u��]���Lj�x.G8��gY *H�ƥ�C��"�qm�>�i�s���Z�x�J$���}�f�m��}e�g�2�z���*�@��F�D�_X��r9��)�	��q�x��B�j\�a�/�f��a҉Z����u�K/�����.'3���=�Q o�Q~��RL�g�;�%'vq���%m!iT��fds���7<�լ�K�*)�,/��'��j��y�"4��M�����Hi��X��)�	}�#'~��1Q��X<.�<�l�gc�9_쇎{N^dY��DC|x��sFk�̠�La;��C�?^���ޞ��'pl�+0¥�ц)o؋e(�I��{D�w[	�{�
]S�A"���̈���x��ۈ
�at���&�q�#�.��Z��F��Nx�K���kX(�-�TSJ������D�BɊ��y��1�@�`vFk�E�ΐ��T�xThC�K@$�Bo����[Sخ��׷_U��� ߉�(�������F��7�͐�>_�G��w���=ste�N0�GtK����߰�``�1��?�+0E�ٖ��rnM���3*��,����3�����>O�J�dj�Y���ƹ�@8�T+��5����So���:~f��A��#W{�V.m��TS��B�KQl��\���Ԯ�+�a�F�I>Du��I��(�K�����|�4C��Vb���J�+'>��2IH�G�UY�+\?t����:�p|�*.���٪����$c�I����J>�h�L���{�2�H�nZf2k�VT�F\���'�1�ᵱ6(���y��}��E����HQ�K(v]�,���ɼ�p�+�
r�q���`�D�S���M�Jm�.��y�٭�x��C6.���L����Ю���1����*�O�y����2�Z�(_��0����E6��T��@>��\���W�����6�B�t]�n�w!	�� �W�;�u	C"��O����
jl�����I��\��L�~�V���\@:�bވU=��RK�G|����{N�̞9K~>�)9f2������|3,��&�&�j���Bl�1Y�����XhP٨�Ch�Tد��^X�C"FY��t��۷^Q*�0�L7r�uB0�X=1RpȖHT�Zn\����85��J� �k���ҧ�[����=�w,�;h���~d� l��s!|x�4��0�P�n�) �M�i��
��Q�A�|��|��.��7Ƨ��n�28�. ۄ8F�����/t�c��b��"�GG~�Ё�GkH!l㈐_���u�#��)�� �G�f�1ׇ�a�5�?��F�j�H당t��9b��ٹ�k��n���;�rt�G�3�A��br�{�8��~ɧ!�;�5ڛQ�u��{qt���	]�p�k�\b��>���$�[�l�8a&�}25$@l����Cb��#�FCxC	NPw{m�B1��W$�"6C?�f;?����4#�R���\C����΍cy;��m����ȳ��'����-�az��0�>NZ��|5�Q"�ro�F_BPX�,�u�e�l�=���P��5T����}K����$�;�ž	o^�c�
�%]��-�RPu�+���$�+���	r��p��S��gUcx�����`打���[��x��X�?n�Psqŏݥ������'tT�s0!?���n~�!�ܐ��D�_<�N��x��Ǻ&G)}��sn��o4��.}F
^���џ?K��O�"�ҒU�
kX_2�����7�.�����GN�!��,�8b���_v�X0\��U��%$_}w���	6ޜ��exk�%���\y���Tx�|���٣1=����~�ű��q�r�j��'�����jTwS�R(+̅�k��^a+G0�����L�e�T�����˚�lp	�޿0i�1/]�>��
Qغ�{��m��o�I\�S�����豏���2��y)� ��{�z��1�a��碑N��|���\7��(EX��"eE�؈�p�O�+�>���m����M�wp�V(r��UIZ���Cn�
����~�ȜɆ$���bj6���fO�j�C������j@���Ֆ���JZ��>�,��7��&�4?�m*B/�f�s���	eLs����|�3i)뺞z8;�ag�j辴�$�Y���@ �≃��=�����[��%+���(����p�������q��2�	��%��ä���wge�� ��D�@'
#�)*)]o�:�E��c����bdB7��U�'Ŋ�t��\cE����ĆYK��D���/p�x��=�B3r@��{�VM�g��k��ݼ�����2�^hJ�M���פq�"y���nƃ�p�~ۅ�������q�}�3�]4NX���|n�ɸ��I�mט�������!ٍˋ�|
@e����,��Q�ו�|=r]w���ҹv_��Y�%Ȉ�C�Zb�{�ꜛ�t��
�J;�{]d��nrT�5�X��s2�'�S��@}��]g����T��ś()�A��Ia� 2�w��nH�r���W�>g��=���a�>��U������٧~,1����?IǮ3'�,�b&KxS�)i����c�S(@��)m���ȧdf��]
"�b�t7PN�2
U�ґ��~�fXo�!��x��XG��K=S
B�8R��h�g"��1(��|1<��PG�m�<�9p���������Kb&+�|ׅ�b�*-t�\y!p���@�&M����wj���|_
����(ͷ�VŪ�?����ȝ2���K2��1�QS|�.k�?\���"�VEjo3p��؄[F3�kxtg�.?&1|�����,]9�ד�ƴ��-�+H����ۚu/��4����.�	#Z����s�UW�bF��8��n��z&J�v:U
f#~��1͗�ـ�0i��9�q�u�RE¼��#=����.��&B36���xB�I���Ӱ5��B���R�=%��C�s���;��E��&Gb�E �7�KДJ��>�++o��0���-6�H�t�&�7��c�'�,5�)���;���Q<c�����^�fGJ�71�snp1��~������-�F��
�D����b	�e��������] �%+Ϭ��wp�a���~U5�Z��֎C:5�K�¦�q�z�����3֣�'��u!y�T��3R��Gy���$���m�����#R	��ҧ1(��?18�iYJ�F�+
��ɴް���d���_�O�ê�Ł�����{{����K7�фJ�4Hpy��$*�M5<��K=6���LW�f<���d�-6�ƀ�9	��]��%H۸�QH��e��#�_c�:���R�	�y��}�~=JPGne7�j�{I�,����X�&�-�nf[�%R��!:���[��ح>����1z��X*}�9�Km��`z��d6W��YA��3wk�uy�t���GO`:܇H`��y,ҦV$,���
��3Iv�Uo�L�t�t0_��Hs֓�lӱ[#R8�?
BX+#J�:W�n�6lnm���* Kk:Pʨ��͒z	sh����9�&��+�(&9�n�i�J�Ŷ�n�3~2-�v�7�͉d��ev���b��/����T�3�ޕ�4�StG$v�%\&w`��}���]D�������;H����(���\�������F�ܱw����{+KF�B�LF3(KH��M�S'u2�ס�~C����lۀ�m>f0/�����׊���t�'.��fK��M2�
��;O����X�9"Ւ��4����.i���s�m�@�?��i{��H-Q����*ζ��3��g~y"����А_�rj��pg��39�:�\ق`:C��m4��0��;� ;qsG���=_կx�|��M�"�#Q��s5��f.W�?��H�R!j^��&����󝮒��Ԣ�|��w%�_�)^�f7״/��>f�+�����LL�yY�1��N6�T��%+ݤ`M�GX�Ժ�7,��"a/���6���~m�e(��ݸ+I���q7ҿ��w�܄f5&��b��3[_n�U���y�g�#SE�ykV�U�.���+���h�8�z��u�%D)�ɓ-V��ϘDvf>��s��d@�q�t?X�+�j�%B����y����
*Z���^0�'����r�VO}z�ǾS�mH1�@����K
G�(��)��8�9�<٬��y��74��: 2�i�4����7P��Ԏ��iG��1k��@]<�8ZRE"��4_u�0�֜ء���ޔ�L�"�R��~���J	��tc���ra���~�EjpH���|An�"+��/U��sY�����ǏP��U�PH�qe�} @��_����]<�Km4_4J4l��T}�/9�u2��;T��FG��E��*��<��E�B���g w ����.7�����u�'�㎾���Q�}��/�	�@}0��j@�'���zON���S�u��
$�|�̛���6��)����'��-���{��)��ia����Ao��MA��)�;,����U�Tٔ
�D4
<��M����.��c���9����&_��N�[�?��ė����X�3��9�g|o=�O���TpW�e�+�|u¯�&,���n;���([�ǻ���"�9���NY�Kf�:+��F ��,�O?U�w��~��l-|�Ng7���`Ŗ��+���Ԗda�W��qB�1�xM�4j��<r��D���WY�k�W���T�D�	�(@�S�+W9ڜ��f��\���ìGx���g� �?_8��D ��՟Y;R�Nbo0���׶�s���1��lT�`�-���ԾP����|/3�9��e�>���'��+Y�:&J����ZrUՓ`�Ei4}�Q;�E���7�����U�|�sA��Xܜ;J3u��"+)F �W��m�V!D�,��ߌu��KP��B���)p��J�B���S\9����p�>�WOC,��3�?��T�s��"T���2@u0ވ�'9/&{FCJ��	�I��t���9�Jj��s���̹��I;�#Y=�FP�L�3����\�j��"\��wn�kᘯɐ�#��p�U:D�!�H�����K%�1(Y,k�& _�Hަ.�q��ڐ�f����=�sB�[t+�1�Z�ԃ�ؔ�-����8�~D|�b��V��6��$�ʝ�~��>��$Q������V����8��LZY�Nk���8����7p(�O3P��k�6�y�U$2�S�����|��}i���Df�y�����{~@�Y�9ZTN� t���у��j�|� ���R/5?�G�I"'���G�,�w K��R��yU�5�ͩ��z�Q���4�.\3��\#�~ǋ�B�Q!�$�ߒ ���$�s�9�iw+����H�&��)�ˎ����lͳa>PP
a���?�EA�%P�r����?��R���mu��➌+E�H�o&-�mRLX��8�F�<9&\������m��L�A־�h������!q��i��XT*��K���"!�&J�H�Qq����~��y��Z�.o=좤���6���,M�.�A�[&��,�~��j�r*~

�-G�u:y��*aX���7�_Su�%Ֆx���2���Ϛ6�\^�`�%�nF�ڱ�i\���Zح�WYKM`�@r�=f�M���>��-/Őbɶ����)���ق�S�YDE��4�� ���U�b�c@�z��u��������m��I�@%��,� � r3�p������'�v"�2�tά�z��lo������ ��nYJ}ї��>zM��E�%*5?�F㪨�Q���Le�Y����mKpL�v�X��h6Xę��>�X�fT����8Q�ϱ1�or�݁m�q���$�����a�����,�(>B&n�`!���.;ó'��������4� �4<~��=HL�_��"�k��0e	ڈ4���#�J0ɤ-�K�bNH��M]����)cf��L�O�I�Y�U=�m8�&��o^�?�
����W5�g�!�' ,f���(��OA��s/*�E��e�1c9��~{�f8A8 /PU�9��OПh����	���[Šd�6�Ĭ�?����ZZԉ?�w�&$@Ź�`"�y'���9Ō�R��z�~jug�uˇ�aSwF�l2yp ���N����O�d2��#FSi�>7]'�ڔMomj�"�t*��|BCt��8����B�Nj��r6Z��X�.�V�ћ��iEB��Y}�
�d��U嬃��򢶡�%�AW�2�,����TM��W�������@�+F�}'@�vG��]v�$#���n���{� U��
Z��j:����L�L��_9I|HO1ķE�N�^��0�cv����'�[�oY`
 �?����kf��P���,����g\�������D$����\��k;|�s'��q� = �,kE�����ȽUy�Ʉ��}��1�7oXC+�6�r�z�ly�Mvd!���g^L>Ә+d�m�G��&�;�W?�͍Y�ß)���/����'�b���*��"C��w��wh�T��)����d�Ick`��� �5�1�T�H)>fs���C��QS��wo���/e��рP0	Ɔ"iq=F
Lv����Ƃ.V(!چB��'#w7�U�ut�%W;��#�kƤ���#�:���Z�J���/��jh�F��7�����E�'�P���%�6���s�ϹK�lV�� +i&�&^�'F��0�p� 9N�n��k;�,�쒜���:�$��V�E�����2�Y���D�g���]�h�� N*j���O��p�����&�4��
��&������WF�\��J�tN퓞[36�b�)��p�^�H�klG�o��=�L#������y&��ˁ��%���,���~���IϫܑD�������{x����jO���,�j	��1<5�V��6Zt������G�)��:�	�����[��'�#s���i_8*��,�g����g�{�:$$�p� u�p���\�L)q��N�(�f��PM��E5��sM٫�P�xm�ECߓT'3�z��
�]pX�l�aO����&�o���?��N��g�Kuޘ���Z�!�3$-~U����<:?�H[��V�?@�����bך������j/��k�T"5�?��
v���uAh�q< ��Lro�+�]���tv��T�T�6T�z1R�������/��~�H�x�䭏��-')�QG��Į`I��|���_��4�ws������-"��(����b����W^��t�@�{p�࠶�
�\�V�2���1{��+����w�����K,:�Q=^��"1Ǖ�~�o�����\�����,1�Wj��ݹ^�q�sw��D0�S�i���F�>���g�i�cJ�65�+���`Z�^+��I4�j���� 5���AVi$Gnp�d�(߇�r��{��t��� �F��Js-wE����(����N�6��a؜a����N:>����>�P�]�!_9�I�h�9)Ľ�S׍#D���ҋ`�/y�b�00,�F
v�#~VԢ�\M��B��N�č'b`�C���)åI������ҙ�(�KL�dЂ����4y��o���q鴌,Ȗ��i���I�zy^e�ɍ�JFb�9t���tC�7����z'����4��7	|{ y�عa钪p9݋�j�v�/�� ��OG��Fոi���JW4É3@ÂIY4��uFH����K|��A܏ur�o�+��hT@Z)~�5o�}A!^�T�h����L�X�Q�m�wF@���>��(ak3�SG����Y�L�#�'nr�wO�j��`vkȼZy�穳�s�j�Qo�e���b����Xf�Ǩ"ޙ$^&lS��:7��R����7�	u��2��ꩠ�f_�Y��DW3H"u���V.ݜO@�T�Eh����Xu�,��H�|;�����d�����1fmm�v��*���%jƇ�2��o5��^=�����.nm�ۡ��(���OF��j��E�^�z�W��9#&|��q�;o�顳o��m�����GD�sn��� PW~Q�>�5<�?^��#�y�1���|�����s����<&��GM=�m)�ˠ��2i��	Z��Ej�+���.Vp����.���h�em愷���{��E����U��k��4��zt�T��Y{�9:��d�����~����<6�� ���`��)���Ѯ��ړL��A(�(GP�	��r��0�����v�j�	к��b�W.����@9C�W�ߪ�Bs
`r'�g���(�={���K>+�-e{���ʒ�`7�\(�?����{���)ݚR�PK�\M4��%я����z=��%;p�ER�]\O���<wfu�IL�I�qӶ"�
�-8�Py�@��ޗd��/����n$�GW8WQ�����ʿ��WE�Yjݔ#R�j��k"�C�[�M�A�m��c�%��"�w@QF%G���XK�~��Nv@�r���y�G�շ��m�|G'ӂ��,ޫ�Y��s �sh��5m��I-���5閲��Aλ��m^�#�����bG+��I��'`��O��`����6�2LW��h��QJ��Qy"�,!1)"�SԴ��ט��j%�k��*9��@֋�W�����ı&`�d5y����$]nG?U�͂��m���S���2 �����?�@�m�|�+��M�5N��GO�����}xjpE�"�P����x�mǋω}���&�y�Wv�Gc�wN�o�������أ@)x}���£�k)_�jʥ��w�h�vtp��MZ�f�ʽ���S8).�,�uՁ�@�*%���lwp T��IE��2��B��NX�	(l�۟��Y�6�척���� ([��A$�o��{<��o�{�J��E����m��l$�~�kK"��r ��&~��x�
���=+�Z.=Y�d�Kn�ᅱ�摃4���A�ҽM��J��_��{�r9�K��?�:6�N��o�wI�h�@��4�z<��NF��.��T,�?�+%��X=���J���!�.l�$����T�������}�K{�ҊJPH �D;:�ȗR+8R������#Z���L�ᨕTiM_���v��Hb��#c'p���J1��r���o[�_
U[D��ݲ)B��9"��v�\g,�$�ž���:���rT�;�A��ևxcz��������`ءWG~���zn����(-,a�Q�F�����(�撩Z�������Sj�$�=t|x���0�uH�	@7��t��;ςx���:1w.�w�j�|�t�Ơ��3�9���St�I��x֛��.8��U6F���a%x�]`w@eJD��U�y��6Id����)lݝ ݠ��#/e�,Z��aת���я^���կm���'{�zJ}1ԫL>O9�m�$�&;σ���Ф�N���}�c��GK�3�Lm�m�( �%@Ja1�ʒ���_�Q���Aݗn��+xL�7+$ơ��_�ZF�m3I���W�}X���1�_C��b3o��������lc�Ӎr��d�,�� �[�p�@w����r���߬�_S	O�Ddd[�=~_���AH� vr����bsv�69����e�α��*����͙ PE|�O������$VU4��i�5y��e7�.\�^�*Z��'MO5��I.�f�ዼ�V�����H�õt�>$��G $��V��qd��Q�n���v�s���A( ���h��n���a5�
����/6�?`��J�i��p�ĝ�����2�B�ᔄ9���c�Z�['��8q�3̳��ZN��G��I���9D��Ulq?=91�s�7�)�W��I��p�"������,�k�kK**�#���q�ЅB��3�������0��[3!�f�V���/)�K��2Dy�Ps��Gֱ��&�2���e -xs��@v�I�k�@��D�B�D��q?R�@⭄I �uޥ���R�Vo��p�a�&���Z��+8��Hc�CEG�����/�E�A��l,��2�/�@��d���ǭ�����{�� �QJ����z�$�4��AQ�I�j4 ˽E�Fw��������s��,f��%�`�����"=�hC7-��G����<k��ʱ���Yh��$Lr�4������9v�Sf	B_�~:T�����9vF|�i���Ԃ�$]M�}`�^>XU�}s�b"���p��%ڗ����X-�[��WY�`HF�]`���-�qa��e�M��c�+�
���V9�P��`m��;����k�W�h������/��@��'�e���0ι���ِ�U�篇��R��>I ��_=��a�����e��ou����\�\ĕ2,qE��*{���?���l7O�mˋ�x�`T�əU?�^ia�J9�߰���M�����a�"3h���y��jjԇ���a�˷����]Î�2��<�,M#`�j�iw�e�mS&�S�J^SD[nz[ �����)��B�z��t�~X/[�:��sx�1��-�aA|������Q�mw&i|z��h;�!&�ř�P��cЏo�3�K_��T�������F�$�!OP���c� ����Q�ѝe��&���Z�@�q���/W�������3���r�>	*4h� ҊU���S ��
��e�K��������C��J�T1^��dD�X ����B�"�����x ��F����/�QB+2���;yaQB<�WX��I�9�i"͢�,J�<�|fh�hFڎϊqU���2��q����Z^�7�ZyAU�lS�z-I�3g���%�"��zd<�*��lq�)���́���
�[܏Fyh���1�f�r�Z9�U��T/+�KҐ���&�C�R�!����ȇf�o���"��l5L�~��)g\���+7�/��j+&�;���S-9���t�-�����ǃ^'}q~rг����/*ʘyC��J']�=��r�V�_�1�
��f���BTڲ���ѿnX�e���^�mw�XjyNMAG~�RÃ���_�����V�ob�6������w⼮�$���B�O�1QYӠ챧l�4.�1����<���&�0����|C�A��t�3�0�K-2l�h�1�W�3�v[, �?�{JW�& ��p`���ABλ�x�b�N������?\:�� DA�
�M��7%�g�ʼ�o�NL2@�6 ��.2>���Pӈ��F�-�|��o\�����Y�,�m ��jAuMP��Y�u��,��m��NW3�/�<���l6�;<���O�9<nw���K����=U,l<�Ĉ.���L���T��'��|�>Z�,���P@��; Eo��V=#P-��l�^�5 �t�v�O�K���xZŻג��A1R�~q^��*��@�����ʓ3XAQ
E+x��B�ն���ܻ8�@�~)�<����K���K���O�t��|Jt������!Q8R(�~R�1'���l���1�>G&�8�Z&aE�G'�q5*A�?:��۳��R�	�*�������������W�6ū���|q�+�4��c���)m
��(�9;�0V9�Q~jᡐ��Bɽ
������,ԧH�Q1+%cr��͛3��jU���{��9���/f�&X\�=�[�� �#�s�\	QU����/{!�CŢK^w�x�+�ԋ�7���h��u�V7ѵ��q0X�M�J�`�e������}�]�J�غj	��HK�������� ��~u��>3��$A�`4�����,�"_ۨ9�,�1>�7:�$�F�2\7��,&����T>��"s��VĴ��L�b,�R�\�K�zA��DY�R8���ѩa8�>�n���1���Fh>"��xSo;��.�������Ë�3y	;$�1O�`Z #ý�>�4fL{y)�_i/z�E���w)��g��֫r7��\� k 2J��*���� ��( ����&�I8�3?O�_m7d4��x�C�i��;V�K����YCm�(��l>���ė�@~��b��Sa�%�H��B@}�J@�(����7���<i��g�沘x�%ղ7Cw���o&�3�X䤪6q��ݾO�L�5��m�|!2R
x=����Z�͹v7J�*��AՕ'����6��MN���H:�;e�ȗq.��B㽰+��L!�����)��"`TDh���W�o���<�n�,��xoՃUn�4���GN�׹�R5窹W6(�����]�r�_�,�:�^5�/ɚY��� b[�~TY������i�R����^G�@k�]/�G Ys|��n�l�L���R����^������޹��MJ�<�qHP�+��-�6_Z�;�c�w�s��=��ivN�{r��|�����h}��sKa�ݓ����o�DS�=O�l���o�u�T&�r�Q/K��B��nj�g�G��܏�ȇ"�yr���ph�����q����_5TX��<єRm|��5���C�@3�[ܲ��]im9*�M�%үv}r�5�!b��!���YK��Nɪo�)���[��X���XHyYa���/��t��K���h ��W��_��e��T׆pg���V:�IޚGdڄO�VN�N0���^����Oal�>�@p�]ِ�G�+
U��ߘ��Q��W��%��.�K�R�f]˛P:�(Ds�{��V�(_�)��&�'l'�ğ���gL�Qayi� S �5��˶]��_�\Tb�N�t@�2��,6�E�y(��H7�N~�NL��&(o�EMd�J�_�R껶�H��0k^��z�gP��e�X�>�6���p��>��/�UD�c�f۞Gm�֘cM�h�� %��$�F�6u�:2�ٕ�Tܭ���[ED��e��vɵ���ț�KuN�I9O5�r�S���c���UV�̜���#��㬷�@�e����Y���vC<q�]��2Jh�L����Ӫi��Ù�`ݍ��2- NlprCn�/����ę�#��ԕ�&%	�a?�Ȫ�ڰغ�F�'Ȼ<2�۝�\&_,u�@���a���؝sΊ={z��
�ZSJ�6�[�Is�
��C�;�L�b�0�(OU uVJ����jZ�I�U6$�L�{p����S9Z��%�Q���~������\�WYY��8 ��������?rC�7T�rzPsq#3$ˤ6�W�D�uVέ�QN"қ@�1������?�������DVCX��r���7=mk�b�Es�˯W�3���>�'�
�`)��Rec0.i+\��/f�4��A��h��r
O�������t�O��&<�Qe4��Ϫ5����X^��H�g4��$�t�@©>9�����r�f�s���Q���Z��qn�Z;uzl��:�`�<K4��y�BN���	���-'��b����c9����&p �1^)���tY���i�;�%�E��{��wFQ��|X�d�qA�������n[��@��$b��f
��G�����
Ql2�����Aݒ��m�d��X�^�� �>�Iʬ�3	��*o�2�O�d��pϮ-��	�R3�/T��I��Ij�Θ���#~�N3|w�0CU�q܇ռi�b���x�*�p�{�h�O�ERs�}9N���4>mn��nQ��F:��a��;�߯5��0��#���J�F~v�d����c�Į�e���- �˜k 8���5�]8��"���[�x�Jw�x5I�Y�{BhbRS�wȌ�|0��x~Ja����lH�ڊ���������1#�*a&�"�$��i
���j�ˢ3�N���!uL��N��h:WMc�;[��m�=腑�|��}Zm���AN7�ܚ��B���������3ozY�d��BG��=���Q�*�ߖK'e����\�{7��i�g������r	N�J�i4�((YM���ݴ�u�>�?�^ȃq�;�`���Ֆ�Ia�uCsX�`8q��j_�������%��},k��MН����4�y����z:ib-�U!:�M 9s4��)j�u6���d.9
6��vx���Y�zD�����"r��pvM�Ø�@դ�/��"�Ѹߙ��f �ƚ'gu����]��}%7�T�+�|�܁H�V�X�}%�;$'G��]��5Ői�2c'j��ViR�Y$/&Xz��4s��I����uX�]Yǀ_�td��E��ʊ�օ���>�T��$�X�k�  �\�a��ӏf�p�����@�2ʾ푱�F.� o�%���Iی��a��#���TQ�<
�V)�����3�g�ut���C0����㬫L�F�`����ztf�F�V6 ��O�nώ���,|&���q�����]��;�<��}u�\Wd�d޺m���N�g-ʺOs���E���>5|�|�h�@Z�����
2�#�83����H���K���S\��y����>�'A#�ñ�}$�Pq�-9���{�=w��*;z���$�SKNx�Z���R�C�%�ė4�!�3��\.W��3��hs�T�;>E2�c5�,���MěQ��d'Fͯb/�K��N[���h(�'*Wx������O��H���S���uFМľ\T��Yu�κ�8��h<K^%3����6�<
��xF�K;��:�~&��L(	��Xzib`���c��9�;�y�b��/��^��T�,oI�a�I�H�k�Ů��-�Z�N7�!�Q<�ނ��|�� �Δ�_�FE�E��"Ox��81<�ca	u莶�F�#�⩮3W�%]��?�e(�@K!�7��g�����E�q��B����h*I7��}�1��
�S�n�q�4�	�ҫ0K�sRI�Dz%��Qş^�A������zW��Z3s���"�ӂb��-��l�W�vP��4d㉟�L�٣z�$,<ة�"�]�$&�#%�8��iS2n��6�=K?*@(�ժ-�{�����|�鲐|/�k�L��"�/�Ax4�3�Q���}.�=��EDнI�7�癆�vV'Lલ�a��Qz.��Q(k}!����zKU�I�#�?[��/Q�."�H�:X�ck=٦� k��<�5����o/����5�������(��ֶoE�f �LH�|@�]r�e*��a�+�h��1�0���^=�n15��6 %A���ۦִ-�ٱB���n�@Uޤ��fd�s!�"L����C֣��aiN�\ ���d�Q26"�1��V�_^G3d=�p�Ǉe��q�W�EC��`0� p���S�H��^{�L]� �u<��Ve�	O_�C3��{%2C��N]jfC��q9�h��{a��u�����U�	T�!���$���i��K͝!N�S�7�TY�B��%���gS	2M����87��F�nyQ�Ü��@J��)#<\r��t��9�5�>���2@D�l0u�������Q��67���[T)I�1k@�a���w3˖[͠*+eёD���̾����p �?",b*�������v2��g��@�&��7���ӣ�0�Տ�v%��eRx>v39v�vWl�Д:��ȇ�R(�sR�@�ʤa�F /	/,�c 4BW���B)gQ���U�zlg ʉ����W�	+X0J��Soɘ��t�fI��Oo~��WǐA���\�x�fU_"2�o*��ؙ�ϙ���;d�`�I�B��.�yPD=q�2;~��⣱ڼ��U|&ƅ9�A��-�[G�8����y�6�5����a2NQ~�~��Ң T��<"zHŹ�Y��:�_a�NNXӊ#9D����K駆3�֗��y���G��9U��b]�����jtH��9m"S��,�@����nx&V��&��*ݯ[��OC,�+�*��&jro���c
qX���Nl+> �>�:���K�n��dE�N�Z�f��	0�(������!~	��b�]^Y�'��Qa���0w��52��񪕄�kr-�Wfh�I!��9��JT+�iva'��`�5��Œ�C�Xq*���[ �Eai��4B�2���uʑi�H���>�z@�O���2�N<����9�h�(Z�����z��^\��b����fu��m<oS�QQO�A.VM��%֔��9��� ��e����=
B@�mi��HW�7o1|>:l�#�!��g��������ql�g"�l�ߟG��}��%WZE
�L�=�4X0��?7W��
9s����Uqd��yW�އ��P��ql��/,(���;DUDZ�<�-�J���[z�W^�d~��O٣ꃏ&�����:e�G(��n�<P��P��,W�(T���/�4�y�K����L�{H�]�s����� hO�W^�,�F~:�a����
6�i,	Q���]g��QP���c1��$/0A����V�����l��t�mӽ죁83v�&Y�ɩ�ha{���X�N��'�F�(���7�1���Hlh�Ꚏzy�z�8M��K��7+��* wL�����R,��x��߾b���=�Rr��2[P̀B}��Qђ#���5��a�c���v�wTNL|������TLp�V-�Z�y�]����R�]�ons�T��|���Q���-/�i1�������j;�����'��LV��ófN����d�����]-u��a�c
�'�ڇ��IE�+��q����{��`�7�����:�,X9�@Q�Y�M��cmw��$;�s�z5{|ӷ�E[t��=���؏�]O�>����\=!�^:RhZZ6�+/���;%��Dϲ��6�����0�N�RQ��I���3���z���61�a���Nƣ^�8�����`W�C�@v�4��[�%Sg�[��i�j�<�Ҥ>���Ȣ֐�s��pZ��J]uH�eH�4T�F�Kn��d��!�����y-�"륙O}#-FN�!G�E)s�/�I0m��:.1[��-)#%W�&ޝ��7��<i#@�-q̙����O�}\^}M��0,|Bf�U���Yf��+�i?7���}�/(�`�NWN�A&'Z`��u$IQ��&�f��.��K�N���5�$
@	q$�#.1��J*�S�x �@�Ӷ�Y6\������P:ۮ~?_��j�[�V�#���o�����|�w݅��"���S ޠ�|u����)��ba+�o�͘g��Sui���?���HШ��)�#�ܮ+������X�9)�**�dr��w�������N�xI�h�
�.�tڿ�S&�G/yCn���,������/
��$��mEQ1�[�z]!%k��K0��i���v�l�`x!��u��+ό����M���zMe�X���9��\�6���x��O�q�lO�p.�!��W��)���Ȓ�2�B�e
�O�)�`~���
�� +�m@rZ���+��v+��z3��~�~A���sk�m"�Z���:�U^@hE��\ĺ���:ʔ#H��;\��2zb1zy=ch�k�ۈ��%c���˂��0!���Qs�Tp���f0x��_�=�����s�&4���O9��VO'h+��J����pt@bh��K��E�%�K�cs[j�1u]xт	����K�_D[�Y(;�6ݍ�++�J��i���(C���^��$Z��s*�ȸ�t�#O4~֏S�h#�H��q�#?3Ql�8����pm�C/;ֿׯ��4ɤ2}o�R'���B�J���2@ߧd�a�/��K�G b�)�-������������{gNj��Z͎�m�T�ȴ<�G����^�6@���<GQ�Z�2���`��ڶ
:�w�V���T2�M�>W�IZ������C#�'NZ*d�
�%��;���@�(�)��Ol#/���5�
3;�<y��C%��S�~=��5k;D�^��<���*G� ��h븽�X���9'�/Q��\;�|� j-����+5����)g�Z� �������)�ڿps�f?�2(�ڥ9y��_���Hwՙ�ae��"���Z�(pg̿��5^���0wԙ��*��@�ڀ�iouC���!��|�D��3�崠�led������3\{�9�aP�2���VÜ<6��\�W������uup��4e�C%	�21���,E��8�?#��[����؁�a��R��t�VX:\˗*��y��9�޴S���,ر�����!]���d#W�x-!R��t;�L_��py��cr�!Aߤ7/Cv�17`��U���R�%���zӻ྄�ޱrF� �M��ˮ*IB��B�vu!d�e}�i��$��$�0��ƒ�E��_="a�:	����x��G��E
���.se�	ʺC{T�>7l/~�*��)!,���}=(�e.��
���8�Cob�z��A�V,朒GSm�{��vh*�]G��5>�P��z���i��ǩ?(��F�"��*�4�g�)K9_�O��Q�Gm�,WM֬��$���I���^r���{Z6l�,Q ��o��!-�o��e)�E�㣻~���X�t��EIB�5���Jg�S��˃��Q���ݟ�C�8�W�kUNI��g0�S��`���;�2�[�ɷ�ٺ3��;����D�2fw����&M�'�z�B�E'2[�	},|�U�V���!�d�L'�'�~�U�U�y�7�I�ӻ�3g<�����!oK��\�M�q��'~g���5ʾn�2{�x�2�#F�g��a�5�E�p��k�e�E/o�j�4��(0u����������ｄ^���_B�&����f⿵��O�4�}�n��4�,v�`�9N��v<�è�M�/d:�"tsF�(ߗ҄����c��K�w���n�+�V\:���y)����y&�k��ͬ�u��x9�o�����0� -�n։�1���^y�c@���'�*!{ O׆��H��(xO���2���}ԑ�yL� ��p��A�p+
��u=��h���!vz,�
=����O���ݘ*�EL�%v���*|��w�?oS�P(�F
ۄ��K�	��'g��1�­8��G񖶚���!{�!�����`w�XE72y��ph���B���M\�f�G��(��[�՚������%{���_9yM\j�������x��u��lR�n�l��z"l�ۼ�#�'�����P�W4�M�� Y����H������z�6�<�/IVkv|T�^t	�7/ML-��l6�]��l���������E�7>���^8�k��e�����t��Ԍ'{)	<�qTBI�L4��{�-L�<�.�fŌ� (7�� +Ce_�ռ_��u��̰I�t���(����i�ti��4����t]���I׷/$�c���!&�%"�"m����&Q�[���_?��BY�4u���b���`��Dc���p���kkQ*�?�EQ�ӯz
�J[g��aG��?��n�V��2�*�� �+���_sE
Q�s��8�@�Dl��[�md��͝��x�UB����o���)��텤l� H��	.��C������<J�C��'r��#�^9C� �,�ֻ=��*)�8 �5I��G����tU �S�X$�\3����ܯG�3btؘS߾���Aa�C�싕��;"&���ޤ0D͒q)���z�<���Ё��պ�n�/�F%��c_�{-�Kk���w�8DO��V��ל�$ �W�'����/�m���̡5��Ф��BJ[�r�5�F'�z�	�<���Q�pT+68���F�YR�Ҕl�ĮoY���T�C��� b,�5b�2j~`r�����}+��U�=��΅툛�J����?��1u�,��`Yqr~!��kYe
.�eirA� d�^V��c9r]y���W��-�3]R���+��J�)��Mh|�H-�����څ+��7SA ��V���֧g�c����������~�O���Ȼ�;��M�#�#b��s��>����X�wě=ʋ<�26~�!�����o0n)��ce�w�L���r�;,Q�1D�2������%n���i }�0���|�Y�4�k�r_z��>ν䤷F�ڻ�ыY�0D���wd�%OQ�Q���B�v��L��;J�p7���]yJJ;Vu�V@�F�,@J�-P�nu��� �&����y|~�˷�1�17�v�	�A�ҴPs�Ӊ���,e��A!Q%���Ɂ�,����݅���k!�*�0���{�:�ְ�Hu����@��65�#-�n=aN��gu���:4�	��+�á�����1��)g��'�����������K�M.N�
�؊�Tg��Ʌⷈ���s���۔���y{�@\�ݸ��2a�Y�� �ɖ��x�b��r=Q�E�[3:�V���p#��-yi���ݲ+�'�����R���D%��c���'sD-m鞼'κ͞+MEO�c]���#�!��u���`�"V�ZSƅ�ᨋ-�;�3|�h�z���CcW��&�3
�M��V��f� ?̔_P�+��O��s�VT�e������5����nnp��E�����Ng���M�|�|�F�Dn �D)��;�Z<�&��T��%�<E��}��wj�"�u�m֖���k��̹�DI����v����d�	�q��%���?��ü+�Y�Ԫ�w�Z6�T/eF:#�i�:I'�L�b���7ߓ�F|O/
kd��u�@;<�O��"�/1 \>�c����-&P�$
�E�&I������������+{�l�ϘX��&W�'�aX���u+����_�E�t�=n�C  ;\���eX�ߒ���c؅9G�0
 p ,�9�,%Kݴ(-��9���p����p� 1<�s�~mBM9��n�7��� �}�Z8e��l��h�\�,���v\�<�i�+A5��צ��ތ�F�i�#�EV[A�������Wwx>��lO��Wm�@<�]gcGn���-C:�2<�O6õ�G�q�J�������r�����C�#�՝�L��"~����5A,��ק�|�����%^���Z���XY��H��*1�/�\���pR�ϟ����6Q�؉���~�
T�u�@\ �?����<����E��v�D�K�&i�1�vh�<�.�)�TR�࿈y�[0��@�J��TC<�=F���&ci�/�s-k�ח{�D���|�I�KU ��� �~����}�g(�Y�1��B\0���ͣ�mBL�_T�@��5m�jRh�9<��EA'o�kLm*��W J�9�����z���'��*q��r� ����sny�	Gp�sɰX�M�ٌ+�SOc�_�����q`%�^�;l��7�4��o%����rFa�+�Q
+�F۔��7����AN����ݡ��p��\L�~.RMd죱�2��f$���uܲT]���m	��<�C~2�ӧ3��/�<x�ǯqy���-oMT����)5<�+�9��O��y�|gҔ�`��v}4�t.C�5�n�r��/Wj��f�ۇ�c������ZH<��nN�q��U��F��9���X����ӟ<�|즇(A� ��f�Q���t;�`�ɖ�H�l����
������?`Nn���4�_$݇��"Sp�A��]k��*X[xn����;���\��\�B�g�#S5�/�&�=�g��QN�36ʨ�����:�����4�W�ǯ|��ނ�u� ��K�J(� ď�;t<�\�1��r�MW��|Ի�c_�#p��7j��� α�Z�ߡ�?�O��<�#��eXC�Mz��.������+��>L�׎�.B5s\�`��d�>�f0J�}��挑�C����T�*!e�P�%����%U@�/�쌱�X;�F��	O�����(��k������{]#׆-g��$|3�������OE>8X)9T�Q����On��SR� �M	�Q\+9�Ev�n�P��L#��?`[�Tb���w����z�Z�u������_��!W:��[�a۾�Y�o�
H�	nh�y��;Vk0ah$����2F�I;
4ѯD�N	_�G#iK�I�B��?�?��G�ŀ���� AST�@�ϑ�:�p	���>��b�+�hr?Op+�-[D�̡����|�b,8�j�yw��S�9 ���I�R��f�Zh)������JWI��G#?"�~"�"t�*����B�mL�y.sWK�T��8�Us��+#���':��փ���5:�`,7�]���F��c�Uf��O"RL V����۰��-B>�䧿����<X��T#ZZ�D��y f�� r"�7�MK����Jo��)�ba�a3��zZl�V��	���s���=>9��y��_w��	������P��1��mt��A"
P�����)w�]Wj͍�?I�x+�t�C-"�Ө�2\�����q��g�5Y�#&*HGs�Ipw�%�|>dQX�A��_]Xi���n��K��.΄��?Ã���x5lW�]7]�^l��h� S�Y"hC�R\7�(���UAS�Ë��z�=�D8��T���8N���s�B�q�L�u�U�8B�cq��[
�BS��䚯�m�F�����[��%T�[M��q��{��࿔�RP=��X�/')�<�Tza�-H�nb�]��X����#|=����CU�_��ْv��W�ߙ��nl��s�Ƶ��žZ��2�ų��>+��2ތ�� �̒�φ��%����T\��;����LW������ֵ"��[V�{P����_� ���<*���c7k~j�o&X�(�͢X#�$�<�%�t���9��_xW��/Si+Uc��N�a���%���M����?����^6ʺ��(�0�WeADb-M��[�k)s"��Z!�~ޛg ɧ䀰�7$�HX� �~��fj�>;/�u]��g ]���JT�����"|�S��M�S��E�b����P��Ɗ�"��}��T�����]��*��4�?�6I�Z�ٛH��f�Gl(�ϠU�"-��a�G�+b�<2n���Dm+i
 �J�?*��oX=�w(ǩ0JD(=,��~�Ϡ�~�o7BX�^C����[.N<�V�Z/_��S���M^r��ֱC5�I�%Ԇ���;�����j�ҥ�A��?�'�4�=�&u\츓5�G���K[�0�::Rj��9������wR�tCZ�#.�wr��_r�b���Z���cNf���I@<Tj������Q"3�D��
9������ Ǡ���"x�	�~q����@�4%��]g�顇���9K�z����ɒ��{4�ǍK��ǋP"���մ����`l���AT%��^��@�D��G��v"s\i��<��r���S��+�c�|�E�T#!;�H;���LW͆s|�{���"=V8�]�Mk�ɶ)!0H�4�zv��bS�F�Xϟ��e�Ϡ��H�U�.�m��g��|�sȞ�ϊ�)뼧��S ��\��A-AF,����Gl�B���k)�`양��d��N��9��;��l�է���"l6�,�4W������"�ɼ��q�b�,���o邵��$�� A���yL�|��O�s�^yu�N�a��'�a����Z����	�k��2��VطN�99�;��-1�W�'�M�R�ٷ��E�p��	��S������)Z��F� �?�%}ga'ķ� �SK��Mt��	Ew91~x��}o��|6
�%�=V��b
l�ﻳ�ڬ��ŭ`����:yPFOZ�.����M���鬼g{^vwn�}oUS&�C��9����.�9B@$�� 
���@��C��`6U�$ٻ'$*M!��'N�_&daua9C#K���;'/c�O^=;b������`4�c3q�S��������кP@��Ƣ
C�3�W���W��_c�n�u�4]���% �9�6_�<�>�
J�R���Z��N���8�1�?<��P%��H�@����g��mH�b�A�\s���[�s�2���[ۏ� �$��6�������5�\6��F��L?�`���لb/kP�A����%怓��I�b���4�V�ʪ���sz��</`9��V��(��B�=nC�=��7▩��v�dW`�@�����T�Ē�%���c�CO73��k�B>$�����I�zO�2E��u��vW����50�'��oY���&���HΌ�r;U�~�m*PF�G�G�P�3�n�:���5T�л�O:X�c�_W�U�g���sspNo�=�����۞�1hh�K�����:(�X|�`�q��|>B���ưKmu�������~��#O?e�D����6�_��c��i�{5���p�'X���S�1sTj+Y;bnI�C3������4���/�E�.�.Q��j ���6�Ht��bk��z�N|&�X��������	�A�~�Tw�	��[4�Jved�=�zʱ"
VN�g$�?nW��i<Q�B<���\1��:i>�)�KU�)�-C�v�F�HQ��?�'�բ�rZ�S7Q�! �K��|�6ޮ)�*a�k���Ͽ�P�k9E���v���$�?�,ws(�`({9>�%���;�ȭTE�N?�5߮}6$WX'���s���"A�Z���@I�fzk��~�巪��ґ���R�|�P��;��̖;��-�����Tr�N�ʷ���(��IoZP�b�^��<Ky��W[I��(2���o��8�	������|��r�C�7ߒ<���q��o�A�I�ACO����ǥ�xN��W=�>K|*�.��>:r[�*�|n����|��6�R�<5�,*�s7�6?7��Bom�l��:�1&e�.��vY}xn��g�VY��=Ǉ�ք@��vܐ��0�զ�R�7�����cI�a� �B�X��5��h˽e�mw2�t�����;>TF���AN�=�Is����R�7f�g�8fc|eI��u&�e�aN�[ae�k�pά!�5��"H�sDܖ�}v���	���A���f-��̗%`����{#�3Nbj�5�.�Wx�N���J���h�&�*.����,}@��NP(%�g�װ�ݒ/�:�:��"�*_h��a��	c2#���������P9���n�۱y��C_E�l�0J����Q���S��(}.:@������N������گ�*Rw\�=��a��ĭ��*��)a�޽<[��i�Dy�Ɂ�C�7�C5ǧ��aWM�z�W4Ti��ef�Г��X�D0�D ����{�u�sV�_`����4��_��H]k��P4�i(�3���=4�CC�%�K��8^HC2m�G[�_X�z�\����C?'[� �w,C�|���鬊>\[C�{d�9��^u��(���`ظ ��oE	�)=�q����,���.`7���!�Ms�(��tC7+���s��8�������(F_(`��NC���x�ˎ��AFV�O��|�qj�����Q��!V����9��%<gt�z��%���4+���E.@��֓�����q�Z�@�&��?B�� ���~�K.�� �{ܱ�E�$!Y��L�����ػ>��@5mLV�t>��Ƕ2�!�lPO�uL�����z�w�x�?9۴�z��k��r���Gv�%�Bc�i8�LKR�ϒt"xjq�D�դ�*�/��Q��<���~ͮ`6oaZֺ�N���t�o]2�1�rؖV��kڒWI�f�������VL��ת�o ݹ��8<���Z2cY�,.��5�ǽ�m~��5�+��Y���!�NL	���+����N�"p��n�N��t�����#��]B�ӑ^�@ǒ�n5�F�T���v���qp�W���!�P5y4�jZ� �X4��1�O�Su�o�B�Hxr�k��do[U��2�Cb�Y�i�+~�A��6�
h��u�v�9V!�mЯ���.����c�b ��w�ΛwjN�:Up���=�ϜHc?�{l�tv�Ȯ�(�:�8���l���������[ެ�H╤k'�#�U;��guc~��C�7�s݂P9��InL�M�]i���eg<��B���:� o]y�^��}�T�e�l�ť�	�F��Kt�T�|�P4���VB�̎�
���n�=��#h�LA�$ؽ�x�'�eQ����4�NRF�N�H���j�ߗW��Cg�LՉ���kDvn�L���ܠ��#�p����=�HA��a�MK'��d*���Vwd=u=�h��O��X�5��Q�[�̪���z�z�䓣�r9��p��s�L���Vu蘿���~��٭��O�
�i)el:�j�5}N�}�����<^��W.��Z�nu?f\l�{��^&J�ͺ�
�g�J��˒��Õm5�IcfD��1@�<2�Au���:'�a�8pW����	���Β�TE��a�֑o�Ӆ`ұ�\#���ف���}�x��q���fw;9�$Ҹd
�q����0
Š7z� ��M�1��aE7��f�h]�eW�:?|]�jT�7�H��9s�����)�(�^��}��ދ�`<�����^Ym����.Ź��[vc���t�{����;�И!@��Ъ__cot���T���R%&n�4oR7g#\�c�a#���qe��åw�[��U���<K�Q�����|����\��F�ŕk8�س_Y8��_�3U=s�r�$!�B:P+>pQ�S��4�
W�Ý��q�'t8aࡒ�C��>�[�o�8���v�D��G�7־BG,jP�I1����{C�zNq��P��PM�d.�y�L�e2Vт0�X��V����ݫ�%dl��������9f��K��(-�5ކ�S���jɪu�Y�`n�Rg���!&p���atY+
l��#�T���muFk0<.)�}Ĥ�^koMp����9X��	�E�NgzWE>h/�q��'%>:ӁD��ʥ�#��HK�Ql����_���a�Ê��=�%�Ƭ�W�(~b	���[�{7X�3���BB�Ad�u�ϒ���W�L�g&��ȓM�t@���8��ݤf΂�"+*bO�`�[�����s<�N�uU��_�<�x^B~ɂ��Y(�57�o����sI!zp1��wl��H�B�J����Ml���
�32Ǔo�(U�{��eH�Ԕ��� ,��Pe(Mڃ�@Oך��鮒�8�ֳA_�>�+v�o�u�%ik�k`���V�Qg��Pў�om��#t��4��7�oC�J�M�)`5����j��rl������<�T��{y�~��X�ձ����|W'��'|V�*�Nx?8����Š�j��L�׺7"�g�d�//��& �/۬*Z�C�X<S���M���{g;rY�E�0xرU�Wͱta��e�:i�*~�ML�͕�e��_�Hj\�|R����,k�ܦIcR��+W}�t+vh��m6N���$}��m���P^�8v=����N�h`<(~����^�C����6��FP��b��`�q��l�B^��S�H�j�B/�&�H���|g�A,��J�	seS�9�)� ��+�X"��H���2S��C\��nJ8�V�x��| 
+������Q�=�`a��}�= g�$�Y�j4��Z���_�k�qFzU�-d���;��MmrK{"嘫��ze/<��P=�@�������ѩ����ڐ5�2��3���_]�c��{Yy�e����@t�yD��/�l礝�Մ�"�ׅu	@C����WZ���@�n�>����9���J�5~1�r6�/�]�x1b��I:���f^�����(��=���XZ��ͨ�xH��CATbd�,��a���5�UV��&3#K�|�4�[�g�M���kL�U�L��'<͟�Isz���Rw�l*�74�X-e�m[wV�n�=ae5���Ň��ow�$��'ş��|Ɨ�S`f���&�͛��ݢ��\����3���������V����s�O��D�Ĳ�wr��3��K]�s�m�������U��x�K#���Pi+���Yfʒ���ULJ}k1~k-�e���5�2h&;ˡ��=C,B5 ���b���3�h�e���? w�bmw�3y@L��7芾�\�k�/7&K�Ea�_���!�r��	�s$�H���B_i1�����2W
� ����������������}��;��h13�[��1����G�3h6^5���`����F�� �KSv�e0z��dE�=��UJC�~��rA�M��A�L-A��]�Y�(�$�&Oƃ[�E���lY��d�X��?��s�� ��J�v5Ή�����DIt�g��������S�E�� l׻k�O��{�9J����d�e@eY��.����yH�����f�d��(�e`�VF)P/�֏�U�O�	��9�$�U@�gC`{�w;ͅ��@��SS���GC����x8R��";��?W��i=$=�kJ�E��/Q��'`X3ݤ�@��Aȿ��vzU�=O6k����V��<���k|��u��4v�ݦ�P�!7c^[�LT�7S�4?;)�嵹U5u��A�ud�B� ���#
E�kv��Qb㊻�|ު��@LPK��Ψ�%���ߔn+w�6���;�p�1��Ț��~�:�j;R{��P���%[�;LkCt�N��p߼��OM6�rby+���w�/L�l}�\9�y9��Z���7�Ҙ7�2���[�7[�I�Pn�㦬�CdH�Cr����� l� �4������IF��zR1�ߩr�������Ɣ,>��Pe.x�DǮ�S����K�	O4w���1�ĉLpF��B��P;����4��9[&Bj�0�`�B�-ޥ������h�0G���z
m��n�R����zj�.[����vz����SA;gԮ� �BgLe�l� M���t'^�jg�S���4C�$5
 _��t!�x	g�%����� ;D5���u�2� m���|�({��1�6~�Y�0���D��.�����0�8k��OOBı�bu��ʧߛWJr&Fq����wJ���O$Nm�n��� ���x4:��r|]E���8yz��� ���)4�uO;�^,M�D�K�0�S�x�5+;�Y/��ǟ`�f��N��0k�Y�{r����
m�0qn�OeXIE�2�O�)�H�'�p���t��Y��� 8L'D��[rʵ�u8n����{/Jzo��=2���kƟn
��� �ˇ��9�ڛ�W�akT�2|��]b��� �x�|�ɯ�g��\CtY9�~�e�DA�����N�hTe��u�p�;y���]�_qd2�]�&)��J�Fƨ��HVb����W�n qCsF��4��v E}'Y]��|K(�у��䥇��!�l�@��㕌>�p�/D�;c_T�q�+�YbԿE�[^_��
����"�O�4> �䁴�6��z�R�ɰ��*��:����q+@V�t�REqY �dϙ��F�9�o���ک-qڈL������> �ŉ6�A�X�,7�}�4�O1ʪ���o�{c����Sk���OX<a�ǥ�6�Όi�0rj���*L�޿����l:�� ����' '�v��3��Rz�4*Ķ�'"�>⟑�x�:�t��[R����$�ǭ7Ac3�LW�e"��~����r��xP�V0��p�>�!��4Y���6�elg��<���GI�ӹS�΁<`�y����J9��j_�I��gy��[�8I�����J"����]*-wT��{ⱴ_sq�m9�f�A+	d�+	$>�W�V�M������ N�b�,�ɏ-��VLݾ�$_�S�Wݢ-�?��=mx�~0t�Ɋ\�fwe��� �QS�I���ߩ�.V�.;R
��pu����ǲk�9pu��������Yޣ]}� -m�7oA�e���q��*
��%v�����l*����`��=��ȟ�kXq��QS�ÄL	|��|�gSv��#�$�-���İ�cM'���Y
��N��0^AT�,h\^��˙U�5XK����ފ�6�ZP����X˦�\�/�ZҦÏ?�	e��(U�?��P���=����]�RX���͢qY2��������}m�����G�z����xj���RXA�L��hm�7�����n]�����|V���ⶪ�y@. �|�e�ɷghB��eZ�Nzi!
�j��/�6~'!������g�����LLd���D��tTT:F*u�X�����{Զ�I�`�����g��Ⴅ�v�щj_�M��`��<sAք���:ˠn�(�����F���$ߣ5�^�Qr�<�ؽ�"L��0B�6ٟ��D�jz�g�@��C��`�Z%>�7,���פ�R-�����!��)���,���08���9�X�9� 2WTl_�tq� ��%�P,`4^�>}s�u'�;i�F\��-����.��9�����j�K+�	�9�ם�׎�X�D ��K�ct�N�?&�@���{�mIa�O߃=7�Ȱs�g�H�=(��(��.�~+��Ġ	���D����-�� M+r+�}����nY�a��#���\$�sxm���6��za��.�ўՔ󁁼b�9�&atS���j��Q��2��U�iਚm���n?)�.$�E�곏�(=�IVE�/��|�^7����2�|?Q��<�ձ	���O~KE��$i��� �-���u�����*Z(�K��"E�!��H���sD�X��>������s��τ�HP+motk$0je��^|Ki��b�|���Y*ч����V(��!YR�W��U��>��4EW25v>,����3����3C���J�>* 8ǿ�����L�9_4]u���`��m��6V����0
��U�ۗ����>9���}��آ����'y�j_Y���_	剖��eg.w�)D�_�i������+"�A�[;��my��:ʵ��-�o?օ���C8����]����=��p�����1�� ����}�\�^O��aw`z�}��F�^tK,;	�>2H����
�RS�INd���TEk���(�s�^���eOv�LC�:֍:Ēb����z���9;��aR�u-�0�4|���a��Ն`PW����\ڄ���T�HK�^I*�uWPLW)��)�̋fI�c�K��_ͺ"�'{qo=�rE ��!�cʞ�	��i@��O����E����O]Ͳ
.�"}�[�����"zU�P���Js������1?�'�Gfj�xQ���f��V�<m��/q���p�v�ݘ��p�:9Ө�QTET�b�����UhFsѪ1�^:�����z�T�N��)��q�����Z�&8����3� �L#&l)�l��lA��0�^x#�D����c��ű��X�sn�����Z���e��h�L�'G~j3Ws�y6�&�)sW���H���������ɠ|v:[^#�����~N����&��!���4�&H�����D��}�I�K�h@A�q����&��*J��T��:���� �"������r������q́=L�d��n�����|�0��a�3#�ȑ��*
� L�{�ޏ]`I*1��� ��c�����Ο&��n]�䪪l�[^�� �T$XWi��-z��ܓ�M�^��7w1���b�h�s����)��s��K��#ݳ�yC& est�(*Xߕ��Kq'�s��=j��1��ƨV�T�\7nj���hD�W���;�zꚩ��RX+��o��ϭ:�nD�s��_;TGt=�k.�U��� ס�lh�a�KPV�*�*-X}�n�p��6d�cJ����%�����c���7���R��i�"��w�t���܉_B��k��o*�"���Ҙd�g�Jg����뉨�A��LӔ���,���.�%�p����N�(���d�gw�2�F���G褏����R	����e��;��"��r�ݝ�¥	�&�t�?�WΉ�� �+����;"�M�k�d�e�;a�K��`��?,��L>���`����
ޑ&�r�2At� �,1��oo�͞����%�)��T}�	�©����MP%F��-h`��țI{JKk	=���ZN�>e��]~�)�O�7lCC>�%OL�]�,ܣO�~}�q+�"�B.�����ɝL��w�Kz�F�×Ő�Їly��V� ��:�Y�D3�^��mR��D����N�)�
n�Bl�K��ߝ���Y��K�1�]F��mz_�aV����E�R _������Q���.o@Ԧ�:s���~*���R;�c,�l�l���T7h���1Yc��Ҳ�����o����f�r�+)�}�b����23@V��}��'ل���0��`/�e���>[��JxC��v�e�'�؝��)޴�Y6`��aa03�0�阶��%�y|��J\�~��[f+N�P�N�d�I5�O����芍��x1�P2����iw��ت`yi�<����I��7wj0�vU��[J�Ղ��3��<��@��3s\^E�2W�(��i�~|�*8���  ��"I�i���h�N�	�Á�?V\�A��;���>|��D�'����B_�,j�%'��wA��dT�;�3v��D�I)O�Y����@�	��,�PϪ�Dl�-U}$�Րn\!(@���;�$��0`�I2���nuZ��hX�Z������*C����S����&x�`�kiN�`���l���Uk�ȶl��)~3���B �67Sݯ\��*z���0@����VГG��w�иö̹! 7�IDt���@\�`ϫ|_3G�5ۼ3�^��Y_��Vy��������S�����E�q�Z䩃�߈�!���WTVsw����7��7U(����#U�� [�y��	o�b��SW�I�2��X��4����
�h��Wn@M�ۀG���gf��L_��WG,��Sx_��l�>:�ővu��R[�c��K#�vqv-D!���f�7 ��f��^C;����y 3�p���t�*���F�8(X��C����-i��*�<wƝe����6~y�D��掅��<e��`�1�9	q�tZ��ڦ�k�\P�b��^��prL�[(㠎#��ž!�_�o9��oB�;xKe�-�z�Φ)�{��L1� j�y���oʒJ�6��"Ta�6�VM̾�z�C(���EEi�A�y	��w7��<�8>7fX�f���(���`AG�����	X�%I2o��AA$>L)�7�ׅ
-J��$��`Y�7yU�q���������"F�)/���d��v$B�� x~ߛj�'i�4T��Um�=����u�؆>�<{�
]޿���J�6:C�; ����S������L�_�W���m�{S9jyי	kޫ:P5��'�s�Y�};T��6����;�Q8
�be��iB��a���#=�d3g�;;�]�F�!S��l7���8����Ek](/���p�7~,# ~T�ӎ��k�C��Z3h�!�?����Be 	�$�VÝ_Ϻ�.m�f���n��y]/j�DV����4����ݽ�`����4�'>c� �ʙ�ީ�J�c�@GO����`�{���	+��������S�;JT��L<!���Kތ�M<W@R{jM�<�N	W��@�m1Xᩙ�;�CS:�@$*�����$T>/�I���=|�g����;��۠�v�|��#?��:=ԴO-�˒1)�����h��,��U�t�<lߵ�����ϳ�T�;�EG  ��>����N7�5r�N��	+/N��fscf|��B�X:쮔���%a@O�&0@�6+[�W'jL�^�苮� ДƟ���x�f���ǎ�^W�������A^����
{�H�$U��\Mkm�_�W�d���M�$��Җ�"�cX��BL����o��������5���������ɩ�671�Dl��]l������|X[�������E�k�V@6Rc�$�N_{��7 
��?��Z�y}�Ek�J*�RѺ����1�b,��8�W\*���r�� 6�Md��M�YCр+�_�-�dM-���I��h��oxKt������AV�͍��莪b��l���ң�WSZW�~�Zٹ�f�(,W��NeR�M�?������t�Y��Ȋ�˸�=�4*N6��g�#Y�����W�zZ�xu6l��\'%�4���53A�q!2����>�8J�cΝ̫���� ~ N�`	����eF�������t�eâ����K�]'7�Mp_и��jnx����r\76��n�cZ�k[0��N�<c�W\�6���z7<��Ϫ�.9r�m�;.!Ѭ�����j�U�~8��
D�S�N`�&U=��m����m��<�x,���x�)1�� %��^����J�P��V����^Tpk���WK��0w�Pq�� ���j	�J��ς �j�;�N�ĞU���'�ʱ��6^����������Jl�*J��h�0	*�3�u�n����J�~_��!4ӧM9�#�_S/B�j)[Ԛs?:�Ts���]�Vl1և�&��[xe��,;����񽫳+ۖlʑ�|r4~��L�p��vŵ�b��(�HJ��:$8N�j8C�ʁ��1H�VM��}�N���u��0��.+�O�#p�;L�@Ii�%d�n��3bUk׼jJ�57����{����jd:ۀlV��,��Rɟ�\�{]�%��eG�杶XBf�2�\߱C��gy��p��?�+^ ���L�rh?A�_>�H���鑅�V���齼�N@L�Ĝl����$���1b�V���NAң�A��Z��#�6h>uU2�b�Z��;�	���i�&�+�T��t��H�!�/���;�:>
�Ϥ�}����9�T����th�����&G��d���3�kVEҧ&;#�qձL2z��~�^\"��&|�wiBAT ��xĈ8�`��c�ܝ&�wF����/�q���3�M������>j�PK|ÿ��9���XU�:�$(	����\��̻&�D��r�1�
�G�FC��B��Nj�+>\-�|�r�{/��<鑺N���A��FߦoRo��(�QV[�7��Z@.O����Q�[6,��N`����V:�G�տ���EG6e�r�CZ�F��Sv#�,�b"�$M�פ���u��ѡ&B?"{ �Yo�k���8?6�̫�0  .~t/1�a���U %N��I2���������H�����M�^��}/�ǩ�Fl1�u��~.\�����@c�]B*6��i1V�<���ל�����k$�r"����ꈜm^�����cog�E{.u�*�V�<%�޵�n��Q��� ��7/@в��(J;8�@(-�f3�m8a�[���zL�$Y��5�P�x<9�_�}�ؠ�-�F���W|���168�fC˜�&;�: �H�;��$-j���h�g����֣-��:G�X&ɊM�k�&�)��='Y�k�DȾ��K��n�lNa�ya$`a��6�/�O�FR� �9��?�}j�r3fAΘ!O��a�	���[u�/�E�9�����<�{ѫ���`�})�����5�s�۶���r���~M��Tc �q�m��|��A��d��X�B�JJ���� ۇ��~�M���$�	�����"$��L��KB�EȐ�����QB�,������p&���{�v3D���� ��T�����6߳�l�Cv������hFk��i�vB]�����k��������@�%i�E��M�|M�i�}�)%)O`�H����� �6�*)�n�����{�(8m�p��{����n���ϞܾX6��TßTQ:ɮb�(���.=�dTr棖��,�+��;q��C�g�Y;RIC��v�_��+Z2~8�N\��6ߛ	+����ۼ�} ��Ko(���Y�PM���6�	��~p�z������5H�m��6s����`A����e��o��Ѡsկۖ��V�����hq��Ob��흈 �ON�.��?���q��ݚ��[�X�NRl�Y4�f"�}Ӻ 1��x���^C��y�ڌ�F�I8��ַB�車>M�M99�*�&(��E�z��䪩�:�/0�ƕ��fw�<�� a:d�ݙ��f-V)��g:fX����܏`���%A�S>P�H�_TfΑc��+i��8o���\hĻ��1�7hp�z �c ���JR���P	=���h�~%���ʦ$4!]/�-_{u_�=��G�ٖ��Ip8��� �M'O�6ڙv�[�6̓��;�ߋ�>#^=y��O�g����t���wd�3��i}e�vO^��y�]%j5�w�`_�j�>��z,}��3���#X��p����%��s�hp*|y��x���E1)D�w����$�_�CO�s%?s���`[/=�xJ\��H�=!�&ocعe��H�e�b��:�'0�`i�1z9/r��cS�Gl��J��?>ehu$;[Q=�p������>��72�(�P���-���H�!��f$�Wo��8�e���V���� y@1����9��4�LCy��L��P���ʱk�(5�3� b$�K#~�2A�R�"��eny�R�� �aL����I���w�E{�p�i]qɈ��n��ʝM��A&�nAw�Zܩ�$	�[��F��FC�vY�P��shm��n��f�W�C,b8zhS��S�R�`�#�G�-ŷp�(�L��2&@B���5�����؂y�d?�q���A��Ea��k\zHL�Qu,ohB���T��*���x'�UzZ��.0S���.��r����z�b�;����ɿ���W�Sm��s�*!�FEK/+wm�U�'���@��,Au/T5N���rI9�XÄwaPAu��]��i�d����H�XvUb���qH|fD�0���X_��!���@U�\_|���k���$���iV�����%�"c;���H۩� ���D4*����뱧����E�.@�~?�{G^��o�-�g<"��B�Xs��� "�嗗�iP��cb>�x}I��@d�U{D@ᅆ��lt��~F�����WO���K��M�\P�o�>�*��YlFַ�*��q|�	���zG̚F��ٌ_��qu�X��f���M��=9�r0t���[�Z0R��/��g�-����w!�!��X�)o�t$���C��@����uR�ޭç�Yߝ�����L��tL�6�7/�/;�)�r�j�(�8�`:��x��i��^U�
q��x��W����9{�bɢ�9OG�c�H� Z��;dl�}��@Vg�*'ws��#)hFC�?���>)Iv07-�J��έz��ˬ�x�e�	��Oq��W��6��G��Y�wd�C�C��|E=��T�"4�� �X����Rˈ
����/f���c�B�u��Bwz��4���_k΃Y6D)Lu��@���:,�=��U�������9[�\�����1����3�6	 ��(��F�{��룡��IqGN5=�u�a?���H1��}�[c�1��,���~�7 9�(	3U��$�g�r�֎`H�ޔ0��&?6���jٻ$q�[�~Z"hs��ۄ���T^��D�͂��b8���7��NCb�����r#��|}cE�<5�S�PU|�E��2�����N6�1N��B��C��27�Ss2i7^�d9C��nT�N��Kh,�	c���}��(��,����F��d�� �ݝ�V&?���QB�'�=q�_L9�M��-l��N�1�)�:DS�j�c�vC��Han�Q���
�ѧ;X��哇�$�&�|��.
����"y�$��c�h6[�M��&Att�4�l
�[�NZ��(�bw��`B��Θ��H!�cy�J{�H����eH���׌������Fi�ƲYS>z4;����Q� �o��ؾ�̛p3nt0��W2�*����CW����ּ��Gk��y@��N���S�����u|~�i�F���Z��}���
��8 �M�?f��G��9l��;��]Z�����0e1��ȿ���Os��9��$��~`��/�{��(2�Ƣ���{��y�seu�����|^æ��nw�?P�4�Ƣ����4���jnܗSCJ�!>��G���u8�*e��l��aJ������n���Qm`uڟ��7��!�u����Zd>�e��j��_�P=����mوL�XX�ң�ܫtq�ޜ��H$u�ۙ����
��&ا=ޓi4fm[y�A!\~3����<�w?�i��~W\�~^���i�N^��3-f%Ȱn��؍���؋�X�7�Ӳ-P�Vg�Y|�� �>�fۊ9� ��R^l��YKT �7p�n�]i���m�`� ��w>�Qn�7�K�G_�Rvl��.�D(�yB�t^<��x��<V�������/�Ȫ��!�6�@�
fGzR4�K ���B{�B�1�T"xA���C�z���iVwsp��I�b@����D�	�psm�s�#KB��9%j���4`�>�g!����ߜ����?��QI=��x8~�B��G�n��R���t��b�@r�K+���ɶV��衽)�G>��LD�`���U�`i�
֙d�ϣ+�`C�u,t���N\w��$��X��U7 H�'�>�P�F?����v��8&����{}�ڎ� ��0 ��O��O�z�}am�>Ө�.kC�X�����?�o�7���a��@Vyg�q5�gL֦��ǩ�q�7�����i���)_�LPH��Yނ#z���C��������@eN�Y�:�~-�����I+!�.o �oʒ+����k1�1/V�Q��u��h����\	?bY׽�һmq&\.tՌ\�Q 14H��o���3xRL|G��֪B���])~�����y�a�8��;8t�/t�e����
��ȩ�IY~&|��ym@>�\
ʳ�9?��J[��NI�j���&�] }s$�ԯB��0�;&�=����.-0O�}.��#-���xf6����a갤ig%~%�.Sq�Bג������u��1]�oC��=Q�E��|���&~�2�RH�τ�E�������r�YiX}d���J���Y��6�3)��<�r��蠌mҊֆN~�P�.�7)�+��l�����$�6 �����J�������rk�+��\�DX���\����~	nb�n=��-S����gÛ>��k�7!7%�����	�KH����t�-�/�#S�S���.��������Tjw�PX1m&�cziy�5*jד�� `xor�bg�[�Y�/�N��/X�|���ōGsmI}�K�}O�$?�>�HŹ-ʆ�d���STu���"���-gUC{�(�K��;[�p4쯒���%EX�X��ZN�����|���D�y94��-����v�-˒�\w�,�9� �z��7�B,s�����3�K$t�Y� dS)���;��J_�tMn�wk�ypz���W�P�Uj�$ p�x��t�n���hJﭱ�
43?�WQƻr��DGӣL�� >�#�@�@&O��y=��o#��Sw@�q���ձícyT�}�3)O�q>=�| �mkG(��h4k����`�:��3.�Y�G����IĢ�>` ���c=�,/d%�����nh���>Esٻ Un��*��P ��Vt�iiW<=IL��H~볞�*�����lLl``�v�d���֣���N-�e��t�6=�-�M馭�e�;A��Vͼr޽9�1��!/�I�&�~���=�Z5D���ϟ��ƭ��x�QDs�~!���#{dr`�V�U���s�f���/{%X���>��-�}���{��T��1�4�No[����V����3�y�W���|
�lL�ٺ�����8�v�����5o�?�x8ϯ>�z~K8�JBi�v���3��893Wq�N�z�`�~�8�A�U'0 U��m����j8�ؘ�?�}��)�?�@M6W��Bue9$]и?��8����6[��5('pg�%�p�#��d��rp�`RF�$��������S������pcgbm��or�I�7E�u�k��>mn�x؂��d��vL��8ؘ)�� �;�V�k+ʉ��e��x:1���RZѕű?9����8��{�T�e����:���C�yB+=���A�/�Ex�^H4.��O�_�7����S���5y^3���^�^�ƛ�'8���sx��D�'_��;�>DmAP
k��濿FLTm�y�]�mp㋱�t?�$��n�Y^�%rE�Q��Z�[ޔ#��@_M.Pzǎ���`ց�)9���*���B�9�-H`��Z8o�5��|ђ&�f]�*!�Z)e�%y��7�f=@	�y]�gԚxۄv��$��!U��$�Ĉ4o|�]E�s�"g�LSub��.�{�ȑN��ղbc=G懺?���E�7�s7P�k�-�!G�b�QX�ǖe��<�лv��j�I�(*������<8B8w&S.�	Q\N�2����K��� i��c�}��Dd��ߪ�wJ���v�Q@�S�_�#v>��+�x_�<�{��5��d3��p2Gx�Z�&H��%&�X Nd<���0�[�@w �O����AK枚��nc{K��6V��.䇷�{�+�~G�n����U6��b�|-���ҕ�8��O#]���M���V}�atb-<��޵\��-��ޠp&��:{��N%��,�-ƕ<nd%�i���e=�����:���g���8��W����=y(2�Z�J$�"��!�7v;�ۡ]�P��yl%�Sh1k��ugI=	E��%�b��\��VΚ��%�H�?y�V}/q�^t"���Jک\,m"O)J�-^�/�L0��X|�&C�|VV&|��b�dՆ�-bYd>��t�<�������فR3�9�-%��WF�5�!|fN�{Z����˺\�g	
)T�9=�;��(If��j�d�B��u���	�F4UB̏��w2˻G��,F��#�{7P'<r��2a��YK�9��߸�!�xR|�H�,��km�.��q5-����T�"Nթ�����=Ꜽ�ܔM�Y�m-Mx\� ��m9Knbc��7ѳ�ù��}D��4Z�n 3���˚��H��WլL����(56�Z����Ü1OQ!��4U�R`sh�����sl���؅��r�W�/�I�4����ݔC�}�/��q��*�� p#��#�����*�g��F�]f$�Ea���I���\���lz2���>��������S�p"-Ÿ���"+�����.�<�' 
�h�3W������4ԉ��=X�0�gx��T�]H]����l�<p	�/ƃ�#h]o���ԋRd����B�i8���� �S���ʦaX@��P�T5(k>��0�L�d���14I���e��<�����Z�m��f�\=ϧqkw��e���Ū$�w��Y@��y��D�ߩ:8�'�-�p�o
[���c�d��r=*kF�.��^�
R�z-,�d�v�nzO�QF��'� ��I�U��T����ݗ���U�X���
%�$�Z�3�b��J�wD`(�$��DǏ���9j#4�!k�n�|��!�-� 5/Ȩ���W��WL����b�졑7��by4"�4"�{���T���&��8iz�^1��B'׷��3������oHp"�;�Ŝ�s?T�R�9���.{�9�J�ުlγ�}e��L��u�n�OXe\������<���9~K�KF�BK�;D�w'��ã�� f�u]qU�#?�G`3��:
"���*~�ll���+��` �|�(��F2d�{�x��N���y5���N��A�g`�vؒ�\�^��u����3�>�oyq��r�x�M��/c�6�mΆ�!J��Bdm=���j��s
3pt�E�j���/Aq0!ƓJ|k+�yu";q`@���چ5��R#m����X�|���ᎈӦ*���4�;"w*0ߠ��`��pE�j�Ȭk��AP2��x��@Oy.���/!~p��N�$h9+��%O���w�b���I��{ܿ%��s,��M��*�&�R�~�/_'�h����Ə�v���|�Ɵ�Ē��
�>��HT�����MI���R������h7�����ZQBa�5gH�F=Tau�^CYCy�G��bc͸��5H�J����m`��S7m�Y{;���.x'�E�0���7+�7w�zv��ݍ5Qq-޶��0w�!�+I�{��pk,��|0E2���?v7(��#�FX�96ع��~��>�<� 
D��^��n����k��&Dvp%jT����g�(CJ�?w ��+\@�6
p�����@���|X�G��M��^��p`�+���a��r��K�oŲ����A $���RA?��t�~X���`[0�^���m,g+���y;��f3�|O����ı��5��R�D��B��<��`��h�2��v�,��:=Ϳ����qc�R������W��1v�Z�cK��,X,��ki��X�4&�>>EȬ���m��.����-S�;�it4ʬgPb��CN��b.� E���8�3"m�@I��q�8�")���Mo�s��}�&��St}�1����7�U�����\8���!����z��eO��o{(I���搐��>���w�x�&�����QV�U�&�=�mZfO��eC/L��p�5����M˚��5�*(w�T�O��B���࿰�'�#<σ�ՂWUIXEjտm��y�=��x_��!〖R5����ŀ$�Ag���P,x���sG�c9�x����'�7֤���+D֧��Փv�\��W`�(r!"�g�O�f8|ɇ����R-��cw���Z�E�>I�&һ�$ְ\��7:��i/r3>��v�Μ�#�	~���N�JF[S���i�H,ǔ�$���ج����'O1qk?���Y�"k��J�m��)�L�^}{�;��]5������&��@5<�=4�J�U�Vq��1�-&Q:8��C�˓<"ȏq��11� ��tO�.GZ*��C����6r|s�Ax'���L�q%=��/ȳ��sE��GsAg����U��%�i�����C#��O��`�s��ʣ���ƙbE��������)���/=Aq*�g"��f�{���5T�U� ���-�8��dF8�^�KZ����zBZ*��D���dߎKg��Y၏@����ym�V�Yq  O/d=)�Ni؄y�������p�bWi[{/?��[�b������V��ҽ�t�nKv���'�7�v�m����CԠ��uQ���c!z�NpNz���e�+��V�J��[��[~�̒P�Ymn��ˮ1ϩ�!�m��tZ�� �U�CM��Y:��Bm�]���a��#V�i6h3�l���-c�Qn�5��69Y~���5%��9�����X2~*�2͐���+��-�쩉�Iޑ���ʷ˷�:�'B�v"�v���
$���"�Į��!����yax�M�P����F]�[00..$�Z��W�I���@sC�Yz�s�	U;#�S%/����65G]�J�S�d��r�i'�� �iP~GKu&�N�i��Aw*4˖ϝ��݉״���߼A��йdSO��0�p�&WXJ�p�f��(9v������s.yF	��|�w��FJ9���d����W��S�	E��	s!a�|�D��8��aoe����J�#�! ����\%�e������#�uG#���J�J:�a]h�� �/n�u{4Q��\NOR��*�:�sd�ʘ8�*E�t~êK9���y��Lo�Z<�#E��Pd:9�E) ���]�;.� =�A��H�_\�i����b��U'	y��f�X۷���W)��b����1�_Է5G�?
�i?��%������t@ҽ�bDȗ�E75�c
ε-ȴ�r���^"e.6!��LV8$��=0������͎���F��Q)iRq��cdzG�"����.�o��.݉))�e�}
�/�f�nb.n�i��Ň�"`v��8����m@e嶺I+s�59,���o�?N������D����
�	#�H�:���-.`č6��.D-��\�7I�Ϭ�g��Ђ9��]� V/�E�r�)$��L�z�`�2N�jA˴I���Ar��靼'��T]2K/tx��B^9:��z���d�o0R�^�*��X��w�A�A���W�g�Ԕ,8�Fs����꾨Ђ�����8�w���L������}-�w^*2Lj��_Q��y�C��ч�.^VV�2��È����.3�,�j�Y�w��	�|�! �^�r0Z��	��rf!����|p"��!'���vt�pYv.��q�f����SLJ#	`b�0[��|�[ϖΞk��l�p���OU&=�p��Ċ����jJz� R{C�%f[����
�^���+�a����� �Գ7o���Fٙ�I�o+�G���P��)���>�y��-z�/)�UsDmg�"p��g��\aI-���:��:J&����?��/���P3�~��r9�t�e��d]�=[A�mV�{eA��P�7�J��t��)_�o4����j��x��]?z#�+L�.l� 5f�"�N�!N*2qt:Ҹ5��6c�V_��C��3�L�ٱҧ�����[<Y�5f��8����)����͚\�1+��b��Ug�1��;!��m�gG�χ�x�d�f��`b9!����oug�dL�l�{�TIR�·�\�=>y2�c����`{�Z��_�J�s�����L��l�!�k�����`G����[��ѫ�ӵ֫�f������hN�%�,_�=/�8�(���0m�t�L��	����C)�:��l&�I��XO	-��� �
����=6���-2&���*% �f��
��bA/RB]�W��R;7�E�,��I�����E�H=g�W���r��� l�����s���}C�l�[��!Όq�#�"K��J��(�j�v*��g	Ɉ�F�M�;0�&�W���=�a��G�b�!���qVM�pʸ8CK���Ow�P:8��;;���	�X�BRgv̈�n� ���o���7���;ͅA5@��[�A�Ju%��b�Is����׵������x�}4@l�,�!:9�sz��y���q �[��Y$��w|G*�*1E�I'�c.�_�G�����*6>`W���W'��8���^z��:`���Պ9>|׿�2@�`׃���WDXn|�u-H���q�Ӎq=����B/�f���ob��[������14�p)�vg�NO̝yom�/6�pX�z�n���]���:$���yf��_�ʹ��Z�ה�k:���$��o�xU U����Iw�8��<������y4�2�^F��嚒�0-�v8�sp,Aѕ�VO�5+�0�[��H�������CU�h^s 8������M�}�_��������GX���ۦ�<9k>�w� �m��]�f�e���+<Ğ|؆�����~���޺��7��
�]�n(�
�x�!ԡ�%n8����	�+}�-n|��4��K~������<􂟍�?=[~�h|!�7�@=�@*�I3 XB�_���9B.ɻ����e��@P�BrXG���y|F{����DK�=�ݩ�HX���=����U1�2�aECΚ���.+���4uH���0��R]0]~�I�&ș�Dṳ]������,�|F����pq?\��,-]6�0bg�v�4��G�d�����~їe���^��p(g������*%o�)��~��R�C� `Z�J���-���v�>$�,��-�O����^�On?�A<��l�<����V��8�i�X2�����R�_���U�&OV�;��?�W�!i)��.�A5ݱ������{�d�>!7l��'N}� 4��G�ڒ'�-�f��cxx�Ua����8�x����q�8Q&��5���I�~�2�yZ�7C�^4���0V����at0���V;wd�uڡ?��Ӭ3���N.$� )��4�-vB�L6�O�S��޺ko��� ����ٜ<�����A��ʘ'�)R��.��D��s�	����XGD�߿�v�U}���>'���#��!���]�^��t�M�i->���"$!ok�J��|�玾�֋-�4g.Dp\#$6E˚�+��Xy5�������͛U������0-����@�e�ݼ��?�GaցWr{��s���Ұ�p�i�Yٲr��S��!\{ɉ��;�xl�=ح�6�����P���n��nm�87���m����3��N�wL[��N�<��9]�Y���Z�:h�OSiAʾ�f��������@4e9��y�o;�)ҹL�w{�F���k.�e@rA��%4-ߚ!+YId�"��6 �]��o�_DC��gE�';iC�>!*5��ku��+��-^@�4�i$����E�b�HI��h���-�k���*����؀C�6�ʖ�6�?zxi&����B��T!��Z/P�]�$�(?�=�KZCDF��OH��L��J^�E��lǷJ7|��lJ�w�XÏ�\4�V�^��Y}�YP E� �|j:��kB@z�Vw��!ұ��h� C�j�j8����A�<��m���	ʢjX�.�g�����!_.���S���2��o;�u^&�EAu����@��J���q 
w�o���0�]4����e1�we$���J�����r���m{j��M!uX�֖�Β��NvYG,�^{a�y�ݙ�YL��^/���"v���Š��B\<3���C��хۑ�1֩��K�~6A���fHJmf����R��#!��C��^o��հ����o̝P�`��d�/4��P�DJ[�pP��)��^��xe�-���Z�k̨oۡG�(�ΛЊ�$ � *�?��8����Ӹ��h_.��VPC 6'Pp��/6�L[���#��d�6U:+��_�&��Gx���ኚkWc)1��?'Yj�VW��KW�;�7f���b��@��#� `�M~P���/�=_M��273�Y�gu���߹wݸ��1�$�],$Y�Q.,͒��*��No����}wy��{��+��8îU�D��0�M1!qgJ0�ހSF�>~[�$O_�V��H!^��F%s�e���q����'���:)6����	��Po�w�)Fs΁�l\�I��ZKo3c��;=�"I��D���כ�E����X�Q+-�]���Ԓ� 	A�&L,��S�Vց�M)����P2�V�Z"��ܭ����������K3�pw��epg�&'�k��D�KΏ{}���Sd�Dkr6-���9r0�2�A�-�/g��;�R+���^� մ�薼#��Z�����>�!�����W	#��n����X�Z�H(�׹�\��wN"\K�c�JEe�6Xc���@�W[tQ/��
��}�
�O7�e�	��5��iU�sU�Z(��ع�y"�!�6,PuI�5�8�z{;��;R+u�s��r�P��~�/M@NƝ�7���.��Y۫æ�X��,��4t8����D>DSSfp�*E�@��X��g�{@Y���x��U�}g��9�������#��U�b@W�g"�4�ψ/�G5PJo���q��?�������^�-��6]�����_-8� zhV���V�K�{��D��V�R׸p]/�
�T�O��_}�F_�j�B�����5LP��Yr޵(�dUSP��Z�/[���B�*钷��;͏�>����Á���=�Y�|�@��0�7����q��#��_�<��N��w�~�k�*��o� �5����C���1��s�`Z���,�����r��^�;�VMy��i�����N?D�`y��Sw��2�ܕ�HC2H�z��E�#��H:�5�>�L ��H�q�U$���g|v�b��n".!����M�9B%؋�b%���7�=8�Sz��!�D���U)�l$�Q(J�h�o+�F-�/��
�KD˹��<)T�sAƪ��z�c��g|4u�C<$��Rm1�ybM���/��E�<�w`�"d���� �E;��ry�6��w�]"�{�X^�O��M�u��yH�nIH��Ǽ�&�S��w=ǁ>�'����cpʺ��Z����/�U�W��·�y��A��.�f�"M�&:A	���iB��:�t{�3�v|��(���Km���W�.�h��i`MĜQV���#焷�)��*3!j|��W�ϭO�9�xk��m��U���ߵ��b6�e���q3���L삅fi?,��4L5��f�mE.�\��qe%��\?t<�J�/"#�ܨ���!_�N��ɇA�˱��<�����8ܣ�$Uw�u:Ks�nJC���T�� ��.��ي�DF8�N��W�*՘�	
x�X.�]�+�i�城px0�/�ƂK��;4���`g�Gp�W�jd�:�Β� �4�h�8�3ry���Z��]Ym������a�K�G��2��?�D3���<���Y���V��B�*��#u1˥�U� �'G�w�sghc\����,�Q�"�W@�1w|���6�&lW����O������ӵp�W�8���iv��pPɤLŠ/�5���d&��7�-o��u/줥�^�")z1O���������r}�6�s.׹ѩeIt_�'�{��&�}�����]N$>p ��ZU���n%H�U�*�ޥ�a�HoU`צ��nh��̕+)���u#mC�q���jZ~�Y�2~�)�h\o�� �3���t�~
56����bk�U�����"�����;����I������k-bC<�����2E
ݺ���ǧ��C�ԛ�4��������t>�]��2c�������4Z���T ������~���+{�T"�]�_� '{������ϻq�bdE
��3�ڝs�p6q0њ!U~�@ƛ���w��z�_�|q�Jj���b��#SC�62;4i��uh�&���L�t���<wR��	(���3��Ľo���(�բIz'���px���}�\���䎺���^8���z{(���a����?;1��8 I:aÍ���Iks�tO��]հ��W�0����4�H�7�j9�}��n�KA��cj-pD����h�q9�f2#+s����Wid?����xd_�t�X��fyqD_�Gw^�8y��j����~C���f郥�׸ͪ�#�g�%6q�
|�4����5�gtZhk^�E�Cڭ��L�_����'f�I��*�W�g��&�Tc��{Qj�Gc�
K̜Q�Bjݔ�ۏ���4ɣ��G�!�ұ���ս�&ױ�� �,S��ʂ]q�;%�"5�}����N�8���.��p%9�q�ˆ/;d�f{Ϣ�O�6�7���6�q����$i~�����\��ܖ?�8�)�jm�I�\%���6�����SfRg�9�)Y�m~m����DG�b �dBЄ������_(*-_=G�^ ,�����֊5��:�P��i��5͕Z����J�� $<.1P�	v����t���A�u�8�.���Q�
�x�~�Q��$�J�L5i2�Vck{�\�O5D�
�V��"�"/ ��p�XM�ѐE�ʿ`Z��"IV!�}ޖ������7�t���L�4�����b��=�':>��#�/�Ŧ�������\��d((!f�Fr�r�I�
a��p�����K/y'qMe���6�s�q�#&�dW���\�\ι� B�;����O�[���5��a��d�7��O�f��G�L�4�Ss�ڑ�وv�P��K��	~F����ۢ���R�x�W#��1;3�(����8�ç�]��P�����ؗ~p2zeg>��7Q����$RK�s���}����w�>k�D��'ru�4�o���H-0��Z�ۍ�jz���9��!��qN�����oc��:,ϗY�:��}'e$�ө�k� 2~�]g�c�F��Ч.m*P��Sx�(
�{�d� GM��������I�����>��3�p;W`J��[L��]���� ��U�	�/�m,���)�O��e�Qb��Ժ6�x확pʲ�d�	�w�b6��p�yJM�.<=�7׎�y�p�3�����fA�?6��D�,j����4� =;]z��[ԇ�,A������a�RJ��@�����V�UR@�ȵ(*��r�¡��b�ĩo8��Q�$: ���$�Ee��n�D�%����c@u}�Q��S�?y���y�;5�WK�7�T�'���x�j���?�ov�F)6��:(�X&���sj2t9�z�GzL��Mi?��[��n�_���ʡ�.��37�ʧ�|XD?)e�1��8������4S@v�_�&��*�����Iv��s��F����V�`_�Lc�d�\�m�����Y�i�(4���
��p���QS��0�E
��_%�v�;i�{Ų�S�>�2v4B�D�èT��h�s�X����h�7������a7��ʉIΉg����p�>� 9�V��X�V��O��	����M����"��"�k5&.N *g3e"���E�V鮬�HQ�8�-#F�3�*�,�B�Ԏ��:�	hp�
+V7����UL�	�}<�6Z�P�3؁��:w�F�U3�ǒ�*\�=��x��u%E�$EYN�Ͼ���;oJ��; �|R��歜�3X����K��E���Zz�VpPL����Ay�D�b��W8u"&S����M/��pZ�B�rƢƱ��WtqõL�w9Ӫ��?�T٩LV/
���<��kEG�S&����\J�z+��w?^D �w%�H�f$�>���X�nk�k!bGn~W?te�GD��6�QCJ�$��>��U>\�z��μ^��w;���`m��H_u�P�1��c��&wn�L���{ZM]�R����_[���)��n����~K��OF��'Za����?�v":U��W%x��z��V�C�Kln3&W���k̵.[���N���Nev��Z��pm�#�� &���}
Rc;� ��E=��)_Ǉz�m��2�Z�^gXl1R%uW}��f��n�1����ϵ0�u	�蓁��WYF�.�ٺN���]�5�P���^\��zt-9��07����Ԟ��	7�^���ߣ�V��*���Lff\�!u�v��>���M�,��x�8i��VgIz'�TD�A��)�1u��z�x8�C��Amh���~��m4�������2��QV�78�N�X�uzM�˒$�HF{mi*�~Ⱦ�6����M�SA�o���#�b{7p�@阍���Kb�]�$������4)f/��K�����!u�Q3o$����Վ��o�ŵ��9����AH����?�d�?�^�����\��3�uQfL�2�n�ϐ8��A{�?�ܽ	����I6y��J���7m���0a�b��1���4j5A���Z6]�1����j�("�M���(�8���r�I��+�,��b�a�:�������ߦ����1ZY�5��A4���*8=۹{���Cy�6�)
�������7�|�%�z��0$r��1� *�%;�d�Z �ۊK�"́2b��I��K��pT��<xϴ�n�㆛��ͽ��*��rY��\.<`�vũ>����w�5�Xy�k���_� �n�����.o���ĵߵ���!�o���:�%A7RS���-`hd�1��#�\
R�/�$t�P�gT�G�6t��7]<��#�����)~�⠨O����kG���X���?P��F�ܺ���i8lr�[�*�ٰ�oC�x2�צ��?騠�'�����r�[�R-Sj3��.U~Oz��Q'��D��h���%��y�����7m�VK����������I&2�"u��Ný�yL�I��Gı����$+[ ?�ʇ��E��U�
C4r;T1ԗ�䙳h�4�h�uЭ� �nP��R�e�K�y�M�-�v�CPX�F�\���pkS��b���ױ:�g��r���]��k� 8�⻿�2�vs�[�}Ke,�ٿ�SD��U|�/a��v�:���i��QWƚZq5~u�7�z�!%'�4�G*��>�����#�r�����L�HOPȯ+Α$Hpo�u���#�7��ٞj�
z��Hu��_8���pu��K#&�L�%���ԒV��iV\T޴�+	�$��/���"�t�5�;qHd��;689��(���0/`@w;�����C��X���8���E��9R��B7e� p0P oQ��g޻������Th�YD-0��Ey�G�?��`�FLӫxْr���N�9?�miJ��a�h���^U��3�i���̋�B=�?�a0��)hd۱h>QM�"fnZVzƬ��m��5^�j�M�V�߼��c{���~i��$Q��> �0�'���e�m{[��Bg�f�v;�x:���8�Kd�o�3����ڹ�:�($S�o]<��� ^��ne��K�-�i���k� ��[:��1�'5Jf�jk�D.��,�?�RT/�)ݠ8�[��"�饀ɣ=�U���[����J4j�&�n(UD[U��}a�fEw��0��7�h���Qh_�bB�Pa9�,�l/��۪��X��m�G�7=������JN�������N�+ai�o�ҥl*j-/foٗ�FF%��=�7��NʌWI�TP���|*E.�zW���{>���K���%wrH����/*k̹�u���<�����Z���l���`�>��g�6i�_�v6��-iXJ���=��h�KZ�M���\	k�åG�Zl�
Ӿ�Ĕ���Ϣ��`CwF�0v�-٨]I皷�H�J�*��h~\�Rj\����(ޫ����d�;f�͒ˣ���˝�Aܒ���ӵ	�b��r������e��c�L����j<9NP*Ϝ���7���W��$�
��)r/¬�"��%E+�����^�۪v�$#
�5��\+�����,�.c6<^0o�����bj���:�@�5�����ƣ�2S��p�Y�z���8	�)S����&0:3�����ԨD���N�8���������7Eo���Bx����;�=M͟P��LƆoh
C�2y�$z�)�1(D����^��x�dI`���=�s������ 9�����͖� ���cHn�y��eK�����w���_����3R�~��@D^��c6eyhF�
�ST�"4�6\Wّ��Q�}�(��MZ
�w�Z�of��b����e������+����ﱺ��k+�?~���S9zL/!���ﱁk"���{���t�������Q������A�m����}��7�0�R: ��<��؆@5fbϒ|qH68cG��07@�F��4��rEg:�U�.��c �o�>����I"�*Iu��,^��f�ю/C��0��s9"��z��]�Qw�g1��*����a�;F�����=1�q�FE�f���m+~-�+�:���0��T0�U8���4��1&ȁ��>W@��t>��Z\θ��l����c_"Q�eA9�K��\�> |�Y��
VS�f�^��b辣y�-����+Z]�=5n>j��v�\|u�c���l-�d�#e*�� ���DP������$@����M2D��y<(6L�wZ�v!��N�{��O���Z��Y5�Fj�J��S�Z	a�E�������I�����5*K�͝�����s2FG�Vy�cA��뚽D��f2�63n���4X楽��� zB#n��4���_80;��?M�Kd�P��F^�h4u�]E��@ίCI`�Q�s/� �V*l�Z9·��\�����߿�ڨV�<5
1yJ��dDx���z56H�A����p�@Į��~x5������{=m�\Z��N3�*#�j1~=(�ڊg�4�����<Z��U''k��Ej�@M��t�`k�Z���׃!8�.^��?�w�|�v<Y��B'�+�@�-�+�_P,LA�����.Z�ϴ�'�p����M�b�����W+�?B5O�|?X�����;zo��B�<��Pົ�y՘9�o��� �݄��_~T/?G}g:ꅁ����-�b�!�)[X3\jR�qġ#N����O1��M]��� �*ά����o�����̳Q�+MyI ^�j��u7MO.x��Zj>˺�\`
���D䪍ܓq\#�˗X���2x��!+V6hp��*��8�&�vȅ7Ft�x<W�����0�j4�ɶV�9 �<su���Z��<�!ۈ�p�Y�dY֦�7�F�Iu�>�<� ��{2�*s\�$���;��"huȵ��d���fq�gܸ������¿�1�5�l7FXQȮYoG򍙮��L�]V⃢Əo���ㄨ��.�����ҵ�d��MEq�%
���3;�:���������-�뛴h�&A!���^�����ފ	�tڥ%����������_kȜ��SEۈBT+M]�k��S�����)��9k �������)���3U�f��Щ�4xi��=W��E��o$D!�.�1���/㫜�_�i���!�Ɯ��׌��	X����˩2f���?��_�%�2��M��j��RN&ǑN�xLKE�Ɨ�~�\u�D\u�0���E�p�xF3a��	���%�z׊�Gci	�*`�DYM���Z~��L�5q�JH5��U��u%�J/���S_K�P��C�dZ��8�u�b%�6���j��u�<V��z���,�Zj$�f*�v,�ʣ�)����)A�.��F�:,���1�.� �H^G�ʲz�Q���|7�˄�^�$��k	��l1=K,�/�  ��[Sv^�3��VM� �������R�6I��I�Q�xYl��9�5��M�~�"�3o5)v~��A�6��S����*�Z�|E�NA���aUۉs�H�@�L���i{Y���W�3�As�����*ñ%�S��*��0�� 5$�t�Ǚ琑�S&�Rև��'�]�~CX���f��z�D
A���]@���B�22�c�z+�-3��`���ba��[D�/p0���$�32�<�W�t����t��*�����JjP���#9���l��՝��M[>�%Gfƺ����l�`��+�~��T������s0�5Ȭ�hbi�r9P�v/_���<y�m��o|�R�w�{�:��/�����	xB�d�,���,"e�Q�
��
�4�J�8�B��#���?8g��yn��� �~,x��}ql��G�Z*&�ag���tƏ=��5��/���X�]����nD��++bDf�u�cF��l��ö_KF$lD���q�/mu��<K�Y��I�Z4����.��.��I��֫�Pz���&���'1-� i�9D�;�|i<�Q��|Ұ2y�G�l~%5��"����k"���V5!���fQ�D�^G_�^^�e���_�x�Ts��:���G{��5Ca`�D� �d��4�����rxd؂�A�D���Ks?�7H�NI� ��>�?T�)s��B��(p�$��)�Aھm� � �掼��U?�-��l0gW0:���K>B���=FN�u;Ԋh�F��)_��(@��:�����n<s�*��]ՙ�IuB~aO~�kH0Ce��������~
�j���v�o���P�NY�tTd(PEBM��"�S+i��R�(8�M��,g(ue~c��!��Yx:ө�����ne-�T��I��LT9i�ׅ#C��.��*��r���1Y]u����S?@���t�^�(K�-	��!ig�I#�pJ���N�J�WS��jϩ�"��WS�E�O��gB
	G		�e�
)�D._�氍���d��m�V/A��Ñs	$�"Y��B%^�A*:�s��b����%P)�(��|U�iv�dc�X����H\��։r�H`�u�ne�ޠ�֥v?��*����J���l�j���T�7��«:֞N!K�NM*���" Y�4�?����dj����!0����|ƩŞ�Sq��ǈI/���P�+6m���pa�`���e`��c�ԣ� ��d�У���?��+�ຶ.�1��q�6b��kQ����!oMs�4�v���)L��%�Ĳ��RZ\5fD���w�I}��֊�'%w��Ί�j�l��A���lm���
��u�ɜ/�Q��C�6��ygt����{%� �:&\[<��<�/b�w�n(�����l��1�O�Wü���`���4@l�klO��֟�w�螾-��
�H���9r/�J	���v�9�/�XF���*�O
������o^���ǟ��ɬ��a ,�z�K�&�/t�����S�\f���|P�<~/&^���~��4g������/ʁ�Bo[�����|5 �Q��Eq)�0lH�>�{�I��(]�V[�Nw�Z �x,p�%Ni�~������l�%���R���Mh�0�h�E,�F�=��E�2b�$Dr�ǥ(�VDм ;��٠�:��K.:�R��a� ���/�p�SQ�s�8}ԃ��sU.<����8� 2�_���NZ�Y�d�lJ�I"�C#�<!{D�kf".���P݅�Zb�6��joڨ)-}�����4�c�b6}���ai����Ȅ͗��L����N�i�>���%0��qj��mE\�|�g���p��$�Χt��������� {��CtA)J��W��48��F����K��m;�(O�@�D���I�U5�Z�O�]DS~.������;������ǅO, O˺d�� �C��=�
������sKq{�&���*���/��mF. Uu0��t;���L��t��r	w�zW~T�~?���7���^ki?ө�Z�U'��跛{�O�I��Ɖ57&�i-���El�nt�uaSr�iӿ,�"���X"��=5�ؙ�ީL����p�%&�[΢�r����ă�2=� ƒ�,�
RB����7�U떩u5~��i,ՄY�<#ZTB�ݠ�xFD�Q������(zޮ9��{�M��	��th���tj�V,�1��D�c�O�����o�����Ln��j��_ �	����)\e>�F��A��$ �����"bKb�N�4!PFkϑ-���G,���&��P�ɸ#˳���t��(�=�ZH���r�M"�ș�n��U}�@��Z� Y3nU%�F��C1z�i�d��;~zԧ7[@�6$�#p�3�}8�.��#�ƾi�z�}\�3dCo�Z�����ݗ�._ܨ�,,��$s�GLe����w��{V�\!��mOT�\d��j6Q��P�3~&�А���#���:&��K�����0�d����8�G��q�T�B������3�Ԏt���hK��۽p��4M6�L���Y�:��-PO*�V�_O(@��Fe�D����\��B��ҏ��v��I������>�yJ����<*$�"3����j!��F��s1�(��yg�(��{8}V�`����³���UaL���؛\��/ڮ�O�z��Jh�X����?Rs5���'܄b[�� pj;�r�l�r����#�#�Y���n�uK����ǿ�3�%����?����/3O�,H����mDh�>QN�t�3W�=*�b�U �\Jr>���x;����*iu|
�5A2.*gVXf�ʍ�^��������Ru��oпh��褱K�I��t$����ٙ��b���+�`Ty���g�F`W��Ln.�!�){}p[U���l0}�cVzU1n��m���5��a�ҟ/���3�٤�����P�Ye�Ǌ 2�U����������4�!�����
+��1�Ǵ'a��U)�%.!���C��K-)��RRw���5=U�y����m�j�*�}��֯�KO�E�iA�/-k�/)'�n�����c{QY�x��F�X�r�)�a�!���Q��G ������A�&G�6�������94�0���=ë�D36.g�f/��z����f�Y8���ɛap|K��i4h
��C/Q��e�Q� �yYf�5e��g�↏����%�kM��ZOm�+%��z�WI��\�%H3�ͩ!�r�\��,)��U,˵:���~��&%��ތ>��r&`ϖ�3�)�˙q�#؋�B�!�e�=s�ӝ��&ܥ�&Z"D&���af]K*F|�
�q�t"&[0v'j*�q�|[_�Q�R~�w=,z���?�+2�/�Śr�����EJNe�;�A���.TI}�)#=g��4E�'�u%�c �E�OҐ��B�T:��� �1��*k�W�㠌*�]g*����G� e�����<�j���:ū����J���>����c�ch���[��=%�|o���	U�d�=.���\cR.�NM�HaK���>R$ɚR�ݣ7�u��t5�i!������eI��n��ʻ�����;:1i�������m-�!RX�Վ��7���N�e�������O�p���/�� ��t<��Ç؊�TӸҺ�_�c޶�ڱ�qO��b�� ��0��p]�� `�x~g�m��RT�9���ӑ#b(fqS�5Xwݙ)/'�3����o�9�{a;R�m���W���P �1��ٵ�z�G}��-!9䕶q���u��)jG�y "EW��A�@�>�gݢm���/2��(��� ,������׻��r�b�+�ɪ�k�Q�>h^ܫ�Kd�.���E���@�@$��'���+e:��SR!�;1������v�Dl��)S7��9�ۆ<9s�z��e~/Ϝ0����Ox<$���g��$Ċ$�=��]�˫��N\�ZHK� >��uV�g�.�<21lyf�8I� ����;��x�o���T�J��}���,���8$PW��N�"��QD�w�U/���J��݈;���`L�Ĭ1ύ �[o�>\2����p��ql���K*���W�S��],l��sѣ??,f���İ��R�_d3��-�J�vG��d0Fǰx&�D����j��� ǻ��)8IZ��@��~��֚G���·���er5��s�=5SWEi(��4�L�R��7�V�=J�^�na��:E�g��rc���S�!��cdZ��{�S�cGҡ�g��4�-�ʅ�p��)}'�Y��$NhO�1�;�h�ɹ�ݶ�P2� hz�&Q�4\x]�Q�G�J�����M��*g��}_N螦zw6"U 
�{�Eb�3�,��<k`q���Pc�H�1B�}��v�3I|��q0�9tQ��`��C����k��	�#���~�2'sp����qb� �g�E:�WL' s�Βd��t�W�jt��������ܬ���6Yq#��A��CKؤS�0JO�]:3n�J�Z�x��o�.�腓!��Ė�{Ls%I&�4�:��{�ћ�	 �@��Mݞ�C��Q�E���/@fX�c[�!7��+U����y[���k�Е��l0kPP��!c1+�ֵӿ̈́�O���\�k[T�kuXУ[Ř���o��sbY5�����c,�F��G�CW��+���(An�3Uu�L��T��N��G8�Pȶ��{��w����ɑ~i')3��uʭ(�g�	u��^+Z��[f�X]H���Z�D�ni,��P@?�ɤALe?�`w�e�}�Ņ� ��$��zDG�U�	5F�*��t�(�Ӽ�u���{�Ϧk���4��/ y׎ ���r��Jد���!e�kYSad���}oc{�c�;�u6����U�̥/�֠u����͜����݀�n�P��&�F��� �����FǨ���k]�@�a�r!��;B�Ӊ���6�&i�=g ё\Efn,@g��t��
��u�%}�� �Ƕ��$���3��+��Ĳ~tO�%��5��6-�E��V�(=R��4��x��Ξ,�і�7D|�Hk�x9X �:ic��.�@hAF�P[����=���&0�g����:�.���i��ʍ˺c]VMO�w�D���U������+�W<�P��G�h׶e��2Z0$���DmG��!K���q�� �®b�{$��O���p\���噺0��"��<mtڇ+��l?�vi�y�B���1U�l�FOlO��5O�$j�nWG�����C�I����'��U �H ����hg[6� @�Z�i���т��:�N���/�v��\ ��ql\xaU�f�,��f�o�[���c����WD�c�Y���OO.؀����
��F�\U�^-C�9.�1�!�j���И��e	p�3YPs�ߤ=zy�p�P�q���X��2q���@P���1��≭�HE���̢����˿tZ��ҒP���1�M��^�!��+,�}���<t.2�+Q T@x�~���j��~�:ŭ�/��L�='�Խ��`&�!��u�
�����B���9��˫
5�J
�-YD��M�����%K���n�V9���_SW=�/��u���p���Di Y׿b�!�H�lx�~U�Q�C�j��U�wr}��ʏ6{b>���3�!C��NoK�z�VE�X�Z�T��L�>b�2��v5r�x-#���/�1��K�y�o�LW��=$����,�6�ǂa�	�eO��8�FF�~JC\�b���>p:"i.��^����n��$��I��0U������!��J���ν��V�'��)r䶍���&�fD`�>߲�=c3�1��\;�a�D�]��:����Y�n�LGr锾?S�,�ӓm�<�7� �4 9�I�c��x�Y[9��k���X��Xɢf���.�>��G�	�q���Ŗ׶z x��̏�>��Xۮ���o�y,�����o�kC��3^����o�|^?���g��:�s�Q�P5i@A�H=��2_��+��(��Z^�K���7���xy�SyqaMq[=��n�U�^T:�:���������Bx�u߽��������Oz�B��9�B���Fn"�ld�������5��~��KdtQ��]3�7��[���-�y���L�t��)����3b �Z�C
X�_���;Ϝg��s�Vh�Q�}�Ȃ@���&��3� �)M�{\�I6��!=R##�(��N=b%��~c@Y ��;��`���'��k���1���Z�"*H�BF;#Xsg�_��:tq��{A��_�l�i��P���4M�oq��wǌ�oR�re��._�o�"���0�Q ��2���H��t����~�G�~�����`��[���W7���������7�����B�����z�w:�7l��'
�9��w���qV�E���8:c$�~^�ׇ8��95	���yuχ<��Ң�:q*��A��-�_��Ϟ��ɉ71�$�N�
��ѠH���
5Lu���,�IS�����eK�#�#��@�Y=+S�%?Ҋ��!�9�Ȥe������>�ˇҨ4=W�ZG��| 2oކ�z0�Wk?9����M?�jcL[��OI��#0ua�2�L~s�xd<EX����b0ϋ�� 8���ҩ�n���Stg{\2p7Q�&Yt���v]�gy<S��Am�F�5fZͣ�F�������t?�.��_0��D��c�[��y{S�gBt]�0��qm�1���]���Iy�9�*�u��D�'ɴ�����6�Sz�=�V���(�&�)�g��<����U���W|��X^��Oi͡$R�P�ܨ�
�*�]Q��[�`�Q����X`�6eݯ�^�Tdz�%8�<���юJ����e05;�}b	�����1d�O��"�aaפ��yB�6#o�=��fKi/&(���O����\6В=Sn'��E��$*3��ĝg9	ה�M? r��JJ�de�T��.\p%4�x�Z�%r���������W2�8���k�˿���@6lzE��L(��{��(q�����~�<������U;ŉr����P}�ڝ~8�� ,��}3���J�bKuv�"=S�Y�yeD�;�>A�l����T&}��P�&LHϤ�P�E2���C�[�� ]狢w���l��ʫ�['ܙ�-�������څ�i!}���I9���\�[^̓\x�F�íre|���+��xY�B�K�y?�)eڬc��+����{~��R(����{�x6�E+�B`@S�.�ed���)�-���"ߚ��Jԣ�X��� ���+��1&��]屭Ԗ-j�Q���1� %�%� ��<Bta��C5�4��+�@"R�s"M��ճ&��T�Ņ3�/G]�rsõiZ�MB<�ʡp zt��:�tT�F��(.�X2�P;��ZYWa�2��o�
��V!����66d�Ǩ��&��2sL8���h���T�'2�,�c� ^��1<Z�C
����m��=��'���*+ֻc���<	��Y��(gY^k����3��oN�2>ٛ��}�I�U����Yӽ*p��r
��r��B��]z75���t
�S���ɴ��e=���p������(E�e�2�mkԁ9��]�$w�{غ����ء��Z�1C�l#�
�D�������b�ǌ�Rl�%M-���`<x��2�o�덁�����E���C�N<��$�ւ�L�����%C��Լ{h�d,D�A�rO��-R��s �]]�݌P�6��߃�	hx��/�GU��ܨ	���"/��Ҳ�;=�79��h,����).d�����U)?9=xy�lIt�]�l*��A�E��m&��֥	��mI��UವE�_��y|.`���?�N��~�T>�չ`nړ�a���l)�a���I�slthN��K�%�l��wBwF�i��_���׮4
��!ܞChS���_(���#�����+["�-�A��T��U�d�spu�2�pq�[RXW��S�lEǁ	�&P}��=���!2�ȓU���&����A��U��P�Rig=EhM˓���un1�>�y��"9���o��y�!�=H�dy����Ռ���br��3�B�Ӓ�8}I�I���P����+5��.z����ȑ���|L ��� �@N,���)ܨ:��:����y��.Ѧ���њ�<Nm��j D�GȘ���DFU�C���C��}��6%y���ƩǷ�`��M�D��Z�"����)-�ո�
��n7^�L�eYP�W/����c5�^#�v7�1s�y��8���g�W���g,�w�Y�#�Eq��(�_����a:�(֮iҡ�ϙ<h�2 ]��5�:�	��χ2V��jİsG󘇢Y�$9ʓ@<��5��V���8m��m0=N_���TrI�u)�0��u�+g�����Ma���?����D��Ng}�APk�.1����O_�"���lj|i�컟%R$_�����u<ix��ek�|��R] >���3!��0���E�1�ɷ�$*��|�����<�(ܞ~�i�H����F���9�S������	����a��?����h��y��ڇ�:��m�!pg�̢URL��_���#1і����ͯP�E�KJ{��s�7ʜ�	%E :��hK|5Ԏ*td�n���<�%[�8j�Df�?�͛�pa�-��YC�uH��>���ܦ-ga���a-ZѱTE�
�L˝���[�a�bW��g�3Vt��O|K�)|�eɝ�����o�	ps���4��Ɠ��;Q�_�#�]����	>$㔡E�pE�m%��G@���Y�Z�,ov���{;D����g�M���|B�`��Ɨ��-'�ԋ�|���VS�a�� W���78W�%�Lէ�@�ey�
��G��al���Ж�bF#���H��i$�/*&�5\�`sC� _:y~�n�yR�c+z�-�-��@�\2+u�=�I���T��0&T�總�[YN�3}�Sd7�O���u�;Ǚ�u��U3�̳�}�u��Z3��ں!���+����n�����'M��bU�*�Q�ʼ�&��7��=1���5��Wh���}ԇ�7��T(���B��_1�g����&�u������h��l�_�5�phW���r����`	6ݤ���S�:8�u��)	��x'	G�]C�r��ζ/��or5$��%7V�nG�h��p}<*;�Bh�M1vAk9���a�m�Δ/Q��弗�@Eِ9�[����!�@$�*F�Q�����$�-�����쨺�a�����|Y����ȝ�ҟ��P�G�_�/6�cDU5�FC��
���G��z��T��-�A�"ܱ�0Yى����)x�`ΝXhh�
�� ��!��e����1�4@∪�$�o����l��̖i|.�WSU�� I�����/�G�����_{�2���#�=]��X����}��q�gq�t)�I�� �ډ��u,���T��eKad�O݅��r���,��G�F@�v�J'���=D
@�l�20x��!�Y� b"��v�'�vir��1����r�ß�=����h|I/��f�k��f�Ǜ%Yp�r[vĘ�4Q�ə-�¿���(/��v�-$�Vw�y�����8qi��9<z�&?�^$�!SI�`3gx�Ab��+�R$�J?�ӌ
������qC^*[,GUo�H�1����]�w@��RQ�ô�7|L�$�f�¸�=I49Vٞ֊=$zO�:�����?l=�q��b^�؆�/1 t�tM^����8����-�i�=�|\D�YZKՐ�c�:p�\�s�6s�����'�P蕴��GJ��g�Y�Q���w�=�e��>���.nfIU���C�ͦe~�dq��70�y���Y��`��s�r�&�E�B2��i��n7b�� H�I���68��5�~h��⺔�k�|*?h3r�z$n$�����N��}׸����M��Rq@�R�z�G%/oI�X��1]EY+@�+h�0G�~��i�^��nhڎn���NzJD@�Փ��T"��t���=���Cʓ.�������F����2�hڴ|+�/mw�WR�QS�Z�k�W�3��|������%�ݹ��ǜ�x���^믤��F�'ʦ�G�H]S�OZ�}^EDȉO*��� �I8uK�pď�y�!l�d2L����pz@JW|�1��H�0���
����E���hL�7�	r<qx,��ݗBO�i��*P5�:. \T�G�2�Ɏ㸾�ӕ?=:�#`�#��NNk�Z��=JCw��І#3�E���"��2��e*s�	[��c���r.nHg�L��vl���#��(��3I���u�lX,~�Κm��}��Ŝ�y��t�nVxTO��Q=�_�<���o���ޓP5�D1o���lu�Td0��]�>k"��`ھ3J�x��e~bi�F��d���"���u�W<�B�4x7����!iz+�B�2C��P��O��߻M����#,d�0h���L�8i�R��kIA{�K�h,�a�#R��J�[�Hi�{�dF �d��֑�5Mq��'�Q�Ǐ�<T�K��?g[Y��Ǐ`��c��΂E�0�O�ra��V�Ma��x���ZsK�qU��m>��h�u(�5R[����I-�	 N�8h.�vϦ1���ô�+�]ʆZ�*{Q9G����$��sn� hU=~#�L�,��6��o4�{��D"����bX�K��W<�O�h1>_����D���2�GP���=�qॡ��XQJ� ܅:�zP<�:EB��A�⳿]Ib�����f�9��]_r%���Z6[�]�H�WiI��Z���>w�~��BΝ�V:F���Rcj-ԋv�r�%l���h���ɒPo e��w��y!K1�1��=��FL�*�:銬�ս�3�%NA���W�����\����d�uAZB:A��Ϸu���kͩ�=����Ջ��<�'�ʐ�js�^'GԂV���Sl	ʊW�e�p�
۵�
���Ǐ���d�r�����3��"I�{��R�6�Ggd�'� �D�Qu�e�D��KF'�^n��b�[1�!*�GI}���ٛZo��Is��g�*�>�0�qII*������ފ��� ^qFV/:4p�wg�/����y �� 9 ''�5�m_�[������u���U_'�;	�Hɸɾ�PW��L�#��{Z�<�p�W�2s����h^#���nD�^*V���h#Ї���m��hY˝v��ټ3�2(@=dR4�͞�w�{���/�R�����!*�fĖ�h�ƃ��sʾS�BE h�z�&Wϟ�tc�_���E�e�F�:��E��>�m�@�c��}9�S[uʯ8������\�R��G{9�&?Y���~F2h�<եUS@J�v��RRѻ�'�ކt�� ��(�@D��j��Q�֐RK��;خm:����\��*ѯ9(���U?*޸�}X`?�OI�`>�T���1�j>]��h@K3r�Hq��j���>=���#�lK21pޫ�G.����
aK�n����uLn�չ�e��1�d7ֺ�b�kp�<X#�b�
{�E������LP�hc��R%�_��e����wV�����4o�N�!j�h��g*K��ZL��p&�9��[=��D��
#�~�2ym���'M��K��������2Ec��ת�yt�����)�;�"��/e��޸��*���D��D�F��p؍0��9�f�a�)�j3�g�̹2�cWv��W�g"�%^�3�Y�����c����s�W}(����;1��4!�_JmU;-���F�ݾ��:J��7��c�Uo��g�X��#�k�O@cG��-�YA'/�N]�>�W?�$�i�w�#���,|�Ȭ�Ʀ'^C ��y�nF��/��Ơ�1E�^��+�؛5%S�7�e�7>��l[Z���{O����Jl ��������R��^�1Ol9����p*X�&����0��)�n�`,�ެ�%��_�;���T���Ǧ��<M�1����}���#�Gr��������St�㳀"��e�C���S&���N�I�)��T�`������Y����45e:�>�sbK�x2d�?�߈����q�����J�B`s2�V;؉�5�kGp7�BXNY�\1G�����-����#�%Z#޴��)�!�^�[�e�J�tG�f;vQx!�N�A7�n��E�OveL���T�,�<b'���!g��ە�����$K�����T�*��-h�������'[�b<^]&��J��9��<��'���٫*��;y�u��lT��"�kBU���7I�'�dh���v��8�v��T��2�����m�N��ah�D_ڟ;R���A�a�X��eG�}�H���z��E�Ϣ��{a=��(6�]��E�;[�i���� $W�jE�Q���l
�Y��I����MТ��Wj�:k/���]�3N�D�-'�G���mY�E�q�����B�҆G������i%U�W�		8�*5���\rX���^{��o�a�ѥ�9��-�(���c�7ɏ�b�,�F��:͇�$����B��Bƺ�$���Ψ�6�ÑB�{W��\�fG�Frh�]d���j��[���%m0�3U���m��fJ��x�}�Mh�cY����-��	�aƖ�VI��"@���/�.x�/l��j:�F�F�/e]r �6ˏ��/��^^�:��"��Z��N&$�����e(>�OM��F�n�S��T�J�Z�`hx�~!�<�wlh����(ϐ��+?���#R*hwME󟡻�-\�mB2�2M��n
�6�nD��gO�:%h�qF�S����	�PuW�����]��]�"�UY󵉘6������1��&�3�#�&H
��Q���/�W��v��oؿhz��M�ʢ�F"�ա���4������TWk,��س�I��"Y��q��um�u�9T����	���Z���ܣ�pN,ib�R94�%p#нZV�zx>��E�_'4�UÈ�J�o���Z���v��ͶX�흹�7��I�j=��͘�-K�B����?�Cx3��4�������� �]B %�ɧ���6�jnNen�t��?���>_���d�I�6����3RL�͆K"���զ4e��ۣ��^��Z?�� �Q�RT�+{ڰu2j���3�`��ɻf�ۍ���~k�F��߁_}C�7��\�g�<";^h�_��io�]�;|߬��"����eI�ʊ#M�d�^y�K�N#���i�B�>-����3�p-^u����+a~�&!�:�02�}�o4�n���ؚeOq��ZS��N:!�oi��[6.�!ڬ7��m��{�a)\��Qk�p͗� Vf�\���d�J���j��+a�~�� ���{)-u%�� V�F���"Vָs��*V>n�i��~�蜗1��kL����R[�XMH�g�W��혉 �>��nGkD��R�3V���f�E?�>7�N�Y�Ca��V[��h�����4��[����U&�<���]�D�����D��ZQ�<�@���)̓iC�3 �y�Ƣ��N�j���=�w,��L��@���e������n���f�uB�4;���y��չ�d�M$�x�o%$�a�C���B� ��g�,%2J�ַ`��Ȅ�2����1�k����=����lՄ��4s� �K ��O/�欱&���2���>�_��|�'�r!>�q�WP<�^�sC�]`ET���~&o�J}g��r��Y`7lYK@_홗� ����j!�P���P�Ό�Y��P>�L�O�r, ����T�"�R�h��{r�8	k���EP���T8�rC�cP�WC��S1>� iUE=r-���J6�M�\,�v�ղ�с��r{:��=
d����k:��s��ц0d����'�c�S9紈V5P'�"XC��m.3w���ӋG��Y�Q���2�0��X�R;/�}��������	�P��[
k���ߨ�[<	x� �fa�.q���eg�} #���ݰ�I��g��!R��Z���y�U 
1�^J�5j֫��P��>��=B�I�؀�	l8�z퍚Ȇ�2ɇ �}�<Q�<��]��@y�l���)�����kd%{Fmk��^�P`h9p�J:�`�	e�u��tk�`��J�i�m����p���o�o��a���u�A��51i�itI����Q� ������2�?ñ"��2_�p5)�b;�DwG�K��da�2�b�\������T�!�q˳b���D�D����tMFoZ�[�� +�zk\�46��ff['�� ə^~��t�\��!�T��q������C*��/��2��e�%5�������9����1�����2m#����q����'��a��1����l�>^��о�����Sɘ��~y-����Z�x`�gk@9��AOi��剭�#=)祺��\�yB'x];���1PT���w�M
j�`�>SȠ��^��}�4�p�����F�zD�������.G���E����l1�a
1�}?�w,��̼�]'�.v��fZ�k]��΁�(2�
]�w'�68�b���`��θNf���?<i3��b�dA��p�A"��� +V����'�z�f2�$����c���1x!@l�+�&vB�l�N]:ƾ� ��� ���z�[����fMܮJ�B���#.P{-j@��Q ��H�uT��I��͈�J��_���N�M��h�q}en�_G�	"��OX9��;t��(�@����]��w7vR;�[S��W��9��$�����Ǭ&�6�>](Aq"�����K�2aّ��f�Ŗ
�y�D�跕(S��kD藶�FN��p���m���id�|t|�E�X��c�[W�g�n�R�Bw%uQ��U���W2�4��6�x���1���k�݌��G��C�n�Z���U�O����<\cDZ���_���O���Kx�e�*!����<�ew*�_{/p	6�O�rc���_�^�n%r�LP3^h��̘/������y��f��GB�R����D�zoǮ��쾖�E���!wl��H�{�1�	7��1��p����K���䦑��+��oq^�%��/����{�ݩ n�{��|u�B�nŲ�ۙ��91��19}J���Y����n����&万��Z�8Q�A�M1�&���b=�	�~ ����hȗc.�1�5�$�C�q���n��aAP#2���n��V�f2���@m�Xխ5�Ound��lP~�����V�0y�ABd*��V-yi�$~��۽A��a�v�F�^�����#YT�g������af90_�ݡ�`��v��c���2��}ګ�'lp+��;ׅU2��ժ�f}�JG&4�����@Ҭ}h�Ur�D���V��DE�_ص��`'ic�f���`�Y�16 u\ t�[�	�<�,��s���rCVTZx�ܝ�l���� ~
Kt�P�¦y�O��O�/�����| ��ru��˽���Q�[/V͙7WLTNU�����m}|1��懦 (
�Վ.&�S��x)D}�'T������&�-�]�KA��3��h񲧉����b3"`r���Q�,l�hH��$
�{�g�R�/{FOl�Vl�Ee�1*Ӊ��<{�py�q&]ƺu�0��Il����aq��%�y�g�p��O���������殝Lf���:�����2�م�QE2�� �����4*N��1dH�(������a��J��2(Tbj�M^��X�{GB�b����+ ���A#&�'O�(rj��}J�V����1|8,�PHnC��$'e0�{��0@ڀ��@<�9wϝzi�|T.ƬZAx��ص�'�Q~�� o'&\&�MX*g-}�*m�	NsE҅�(M�������0�>�l���8�nj�G�+�,~H>���xVP�bLoP���E�����{�f*��1ǩʏ�m9N�V5���D����hg6�پ��6OP��fK9ypя[F�c�趵U�|W��ԁƯ���2����"��7#��_؇��ç��٪#&'X��@��Gu�����MDMqx�2�R���Xk-;��n@�f*�]�Z�N�ۏl<]4�t��VU�L����B�
��>������Ob����q�~�M�K!�~���]!Z�h�9�/���ܽ[�j�A� ���;��\�U��-��J¨W��g��D)�.q�e~HU./#�X��	�{iꦢ����-#��p�s�8�v�zZs�3��I��μ>9|@�4��x��k��`�ZXd����\������i ��_�ݷh)�y܂s���4�E�Vz�b
��޷"U��]��ld�~���k)(��H8�F;z~�)+Jg�܇"?@���*K6�D�c��@�t�_�swEk�7��oDi�p���E�����ߢ�:7��4�c����g`���D3��ѷ���QT�Y)�sbe�Siz�+��〦gZ]�]K����L}Ed���k9W�Z��D����y���U��Oa
`��|�g�=s��������G�;@�*�e��2T?a�6{���b���7� ���A[ժw����}������q%/���vd1�q.i��=�5�vP�{T�ui?������D���}
�GJw�E����"�A_80f�	^�C��e�۳�/���9S�:����h�+_,��������=D���TY����ii�ޘl)=�*�)���g���V�mZ��A�6��G{��������]Y�}�׷�]9�ҩ�jO=�KkvC�<j-��f�Q{=\�J<6v<�<*�G��
��:�1;�8$E6�ǧHT�!8��
wz��k�y�-���&Ƹ˲���K�^���/���Y}��1j��Ƒ�4��l
�'���ROM	]ӛl)�zr8�oڑ�E._h'G�%�}��ɮا�L�͙�����P^��CX`��Vz3�#z�<��k�#Oؽ_DF�����<$�C��]�n�s��V1�dg���έb�ܴWB2�T^(�h�¶[M���Wp�/��a{�T��r����=�޳��*	��W��D�[ߪ�����c�$��G,�;�е�xf�u��\4�#ǻyӟ~���6m�/��ډ��y�&V�M��� ��؁	cvu�Ϻy1e-(\Q��%wv$��6��tk�\���'�$+�y���1�	�����	�=�@Ԧ~�v(��!���P�uwVO'@�� ��٩��n!QT7h!����v�了�����2�e�k�7��p����ȼ��b�<�h�c���P�!�����N���'��E/+]Z����V�J�ƽ�L�N&������c}��9��Ym� �A��������'jd^g]���*��8��,�_��P;�zVzF� ��_^1��c�&'��L�vW%�G���ԉ�C���d�o��ˢ9�٧#�������}���)�u�*+S��@}�����;[P�af��	|d�C�F�ֽ�-Mu����bM�xR�W������%r 5 ��$��OeI��4��[��ݧR�!�)+�"����$pό�p�5ߔg�
S#V�J�/,w���5�Gހv��yQ>���,�v���h_|Q��<� ��c�4������<��'t��ڞp,��n�
�`����A�΍�L��%m��<���\��G�j�4�t?�f�λ�|ߦ���(`�/��h|h��B\�o�<	����y���6Z�pEk�p`�<s��܊�����V|�k���`F�ɆS�M�d�HՖk~��u���n��H��`4���i` P|�]�':�A|x&�@M47#fBji�r�k(��M'*L;u�u�WΝЍ-�Z�`�1������+�0�[T}t�y�R�)���9�˄+����/~�����:<�Q�T��Kk<x7��#ӎ���aKq����������sB�����qng��z�e��n� �da.~�@�o�쟠G��n)� ��LT�K��3�5q+�A�'�_�hŏ�q2�bHN8i�=<tn�X0D{r�JSR�������܇��pkt��<})H�u��{^����'}z�K����Ğ��?��d
.���'{h;�R�Ղؗ�R�P�ՠ��V� Y�7��8~
�9(w�<��N��<9���:�D�O�O�x/�V�L��6�6L;���t�:0�Żp��pqX�u�s��5��H�y~����0����Ś=Y��Qg�vӒXd\��a4gd�!ь���@h'o����i�Ju��c�՚�5�fKVc]v^���-I<�>d~�+�p_ ��M� �,D1q��9 -f���3�t ����#�B�{��L>��3������,�����y�O&Kܱ��Lh�I��!��Ȍ$¨^�2o�̣Ի���:�,M��U"�/D�J�v����f���1Z�'Q{/y�P�&�oڄi�5�_E�Y{{>���<��B_��/�9|���JF_������#q��ZQ��E��g�&����������wl]ij?S(�:�"�a�أLW�Q�,�!F�^�S�����	��+�S%7�,M��W��)ԄD@u+.F���麁Ю���8'���n.}�ۋ�L�w��7�,N��;�!�>��y��}���+��Cv�΅ںѵ��2U2����"A��ʁ����I��T�/i�=��H�V�(�uޘ���~�'�Ѱ��.�ڜ�� ���
��G�Z1����S�_x���K��Ϙ���DV��1��f�X�3����C#i�l�0��k�3�||����( F�@[;�oQ��ȉ�����y�R*�����~~w^[|J�MT97#Ґ�x���و��K�)r��a�Z�3�Ls%W�X_��g�O
�hK�)�Oj3�A����3�B�a�;��}A��/7bf�"Ȫ���C['C�Xb�]ft�<Έ(q�WF�ʕ�sό�oɂE� >���
C�q�SW����ewq��^�ui�����&�j_�ĕKb��=��W-S*H��L3;>X��*�����
$�O���wl�o=��F�����=�����-C��v%ې-L@��~p�օ^\��Ѯ͑��d8f����:��{�8��T�p����sVdt��y "E�IsA�VBG�VQ�����^\��b�t����3���ױKUE�a��}n#YN�7�	�&,9U����B5���*ҎE������K���D<�z^����{$S�-b�u��l
�������e��ڸ�##��|=^���[tƭ����%M��Nݨ�F�)Ԛ��%�$�{��C��8�mI�����Fu�wsR���I��s��s�/��ұ�w ���<�k�����	>��%6�v�B\V�����7tN�p��54���ǛK=g��F��	�ˍ�
B�y-���1�n0^[r�$�VJ��$ڐ��wfk8P��M��B�ܓ��B�=����e���)$��KEHn�6@�C����x�u�}�(<�K8n��[�E�:��)�\	��f3��U�l{�m˥�h��e	<h��iWI����6�[>�#�9��BΞo|�'&��0�k������BV�/]*�V|MPs��̏��R.0%T�j־Qu�
?�'I�ő�0� z_Z͖�ܪojHϕ���,�g����������w�����ܧKX۸�W�\����2���G��0qc�ɤs��	�Y��f�P�>���v���A�&���q�^��0�N�ȑ�{��-�J>O���>�,)B���Q�?dq��Y+���^(�^�΄;�4�<���)����!|��ް�界L�6/��
�k����Ֆ�C���Pb�Gr4'�wN I��f�=����}���;C�.�l�6��� ��/�E�m���YCA��Ν��H=Z��EL3�#�E%����^����_%"e���	 &ҮA�_������8&��lr��#>�k8=��Я7pc�2��	 /=���do\�^ZÌY�DU��菉���G�v�RLn�|�.���~��ڂ�XYP��r{���Up���(< obA���d�5����d%�8���J]����z��$Kv�Uj�҅�5�gWPݮ|��U�A^a�/���[��I�,d�T׋4�����\gfT����ZRO$�f@���O"�6�s�kQ�-r�ȑ�����c[�)�S������u�oF��
m�N��3��^������"$#j�`\
�b�%u�*���8��F�V�0��}�(��
�6���6F}y�H��FNZ�#�����j`�"eN�֔$n�KJ�n��:ٶDwb,GsHPR������n'*��>�����Rc��<@o3U�d&�$4"�܁�:yЉ��ԫу%�%��,��=zMy1�� dƝ�Tyķ�������1�9{R��p{5BE�^@W�&E�[[��#�=���[����9^�h��̍©��h�oH�|7valO	�C��9NE�v�.qk������~:s��\v�������1��� E
�PisB�V��;�B<t�K��s��Q��]�m��D"����m���v�8��l,_����S���q���S����|L�B�Z�)��k�UlQ��)�����x2"~���K^/u�ػ�R*�8����Q-���K�>.���GT���2�bl�Uj��I1�1��8��|J�c6��m0�����B�}N�L)��?�m��҇��+��D3�*�J��a�:`�)�lO���k��������O�P�7���E���cr��D�c8�Dm��.�aӱ��&ug��A�k��f��\�IK�y�Em�T)*6��W5_S���)�QX�O�?!v���� m1�6 K��&���4)[���CU
K�z����#\9b�^Tmo���}n���I��=D�h��qr*[�"��g�O�X�=�i��>��V�}{B&���Jx�a }��9��{��N��h,2H�İOcv�����h���&��Q�穓�՚�|9S$8^x���G���҂��-"�ߜ��Z��ʥ�\쉼|����q�S����P�����P!o��o��3`&��_�"4Gڪ��>]���B7���dҟUb��H��M�DS�}�+�8���H*	"���\��P����#@�x�`�(6��{8�l��ae�y�����r�&k���h/m���"#Y1#.��;����w%?wlO�R�2�Y©*��i���](^�1��<4���}�Y���n0L�����G ��O�X޲)��g� bJ*luI�#�~�m!�<�����
�� x�xAg?�Vw�kѝwf������ف#��	�i#�:z����L����M��ӷ��7.@���L��O�4�z�2
1:Fz�CK��/�!�F#3��H@�|4@��&U�.��!�/~����"X���ԋ�TK�:l;%{87��EM�"�8�Q;�� ���;%_x`����h��9.���4y�����m�0�JyWo���	ެw���P�~��~�_/�Ɯ��W0h�͊��< �Z����,ye�[�`��D�~�e����<=�Փ�G����J��@,�#�� .���9Rupc�\��Lq0"� �]�o�Ӽ־��hk���5�K��"��ѩ؎�eJH��R�5���Jo�QY����>$�
p��j[��1���3 �=W�\���Y���/x�P�(��dы!s�"|� 	�_�`s_������,t�����~����9��SK�	X�(v�ۄ�x�c�fXC��zb]�ߐ�%�|�M;��$i�O���g����X�B���A�w�w�[#�h S��a������4	�~K7!�)�A;���x���+#m��
U�u�&e�*<�]~�A5�_���>�����������fCF
OD�W�Uͧ�3I,�$���J���LA����ߡp{����������s�1jʅM9Y�kB^��]�[�O�Z��̧ن�V��I��q��
��?��4[4�����)X+�̣~����9H �K?��%�e�N��wp��R���I�4!\����*@:�Vi@�[s;�r�v�
J�#�%P�F��7_�uE(�kI�}D?ױ�B��������t�n�&C]���Y����}=\�#�}��Yx���k�5�*��}Jj�x.�)ji4ԉ�'k�&�ˈ����	��¹������E����5���X쨮,�1�FY�gF�3c8�)�*�ny�;�/'![�r�t l	��]P���C���5��>�FO�x\BaJ��3�v�Fw���x�9��}Yρ~�o��?�\Dn%���<��H餮�����	3 R
g�b6�9�"�c
B�����vU��̪��Lk�1�NT[ލ��d��G���i?���7��i3��ӣD�?M���1+�!�]�LsZN�?ec���!���|�֛8Ԩۉ���Xc|	���"͸�`��o���ޗ�Ϡ����t#�!�Ы���-�Ž_�����-��yK�;�|��
֫q>��~�hE�P	E��� ���F��@��
��bƬP�/p����t��U�A��t�;���1�������V��g+�ŝ���+v&2A
�0�H��v�Dݲo�wz�!�X��֔��O|���ԯ��/�4�n�[�	�S����}�#�`���nN�Pк��%�c��K!��^�*z�LW���z$*]�+㻖39�"Q�x�}���._To�Y�_pM�t$&u�"�\�-�UjV[�f6��=F���]ZD��y����3��>�Y-���OKe��.�B^=��_�G��ڒ%����Q�f`���|�}�� �/��E.�-��� k�}���H�@r��'�6�5�?�x��L�|��{/�E�=��q��]Ӣv<Y*��1�X�	�S�!�9�Q
Zh�����8O�	���������!q���y��:��A�UJ�R������w�9X���*?;����M�����A�+jsyI�����Egء������c}�����p��_XMMzx��v�x�o��?H]i����J�2K߭e��
�H�ďʯ������.`�`��J������0���E�-S���RT#M�nk��9 ��$��]�4^�D;/f��K,�>].�x�L�<�����X0WO{�3Wf��j��ì���I�����.��@�k0\-�H-,@��I�$~d�>I��=f@K�UԦ�y��7�2a������C�SQ� ����A�I�� ��W,�+��DѦ�b�ض�Ǖ_0�����	������$-��ѿ���^mt������ԵGиp��G�x��
���%�z Hw�0ȰJ���ܖ{H|@���;�9H꟪.���� ��x��4#�A��W-�lI�+�e����ҒB=���dK�(`0W6�!�|�r��h<�%^�tp�fY̥B��'�A�4�W�Hᩞ��NeC�S��H��"�74U��&[��xtގ����A�K��Bw��c�΀ګ(�QH���(d�D7v�"�/�v^��K��{���y!�2D���+&HNn߶4#��Gi��^�wv���ܕƱ�t��/�s\,�T��� �_sq	���$��+�<qO�ֳ#9�&?��6�����������	�+A#sPj�&
�R ¡���+��[��u@��G�`� m����|9�J �d�6��Fd���B���ye�Wtr1-[�Z�P�1z�[��Nf��c��3��Ax�t֯�^������󷳀�����Ϳ'p)����j�3����7�.�.��7!� 6~�ǔLU�(=��#��$���ܻx��֢�S1��,�y���M^�=�me�#�U��n�C��s�A4tV��b� �:��1�9�j����;Ŵ�=�0h��va@�}�ƺ1^�˵	��&���p�%*�ֵ�q�3�`2m�����Hc��i�=TnK�a��ǂuj���E}��A��d`�="��P�z�d>P5a���w��=4k	H,˅���S�&����Y�_�[z�U�W˺���Q�ln����aZ�����!�>ߩf�o�շp�s��հ AKA�r>��/�n�y΁_��i6�����J��V<��/d��aK���x]��|N�$=��Vc���/,ꎌ�׶�V� ��t�gG�Fc�t�o��q�5�ٔSJ��[����Z�@��=U�4�������048A0a�p����=UU�t��U��׍�Ԗ�8��e���A�W+nI��wݿ������*��hu�������~�Λ[`B���v iHU+4W�1k��<��-��]��h�H�)�J�$k �,DZ�oW$�s�!�9��=��9M	�P�Ka�m���ޑB9G�jȑ�2m��߼� {���ϼ{'�f&*�ki!Ex��?���x_���xrK�_m].�o�!�N^K]���:��N���byD�M��x���ǩs��y+z�}t���ab��i��ϵt��=����;��ꥸ5�����;H�+����%qg�#h��G �v���j,v�"'z�j��d5��d,�3H9<�%�]���z�t�����Z�&�g���1 ���آ��7R^^ n�;���q��PK_�.V�I�Z���U>�@9d�u�s�P3<q�|��g~l ��O����%�ɜ���:� W i8��%_�e��4
Ah��F&��/�O��tp|gzݐmv�@��i& )6m���<�`�zZg�o��=�ؿ}��e76�H`m���6ش����y	l�KEՎ���w~�8<�����j_��k��yxm9<�mý.d�rt4��-T�6�f����ew��Ӯ�w�SsP ���11��AiE��O�ym�A���n9Q@ .u�%��Jn �)] ��D�<�<����b�R� ���[�ڸ:����ؘ��Y������ܙ!�@�SA>rFC� �c)ַ<�
Ϛ�_�$d�h�"O�Ŀ9�}�-�XH�yH��:���S u�C0��L"|�#�SV k���oϰ*1<m���]�GJ�+;�������%+.%�/O��8���~'.yC|&c¬Vs�͓�.�`���S����R�<"���ǥ��b*������������.�RZ�;$�Y���F�p��A���H�#��s��e������Г5<�����r�i5ա��7Z}���g�Ң�Pty��g����-�a�g��u���EޙnspeV��J���&UE�Ը�[��/zM`��}C�1NV uq{��E��aY�|�Y
RH��>TMSTx���C} @xGܧ�A��i�>-N5��Y�0���P�Z�L�DA7���L7�*�B��?�~?!�G�?Y��g��p'R����t	В��jE�L��rX��3����l��@vE��ɏRHQܟ�E��n���B�'���6Jr
�_�b���<���!����mӮ�X��Ao#ř��ӣ����+��b�\��I����Nc�8'BY�Ciy�6�W�T���ĩ�U	
���Ô��LbΞ�v��Q���Wa~1�%����3IHZ��l��8�� Iq�,����'v�y56le�z̤����-�(�� 3�B]ini�A�o;F����<4��m�	�cLNh Ymt�cfr�@��X�ep����*|O� 1n�������ݼ� RV����(%�g�_��/�m��7�Z���e���b�+,M���Ad��L|��Zr[�� Z�`%�}��fM1+���5�A�/������Wt���5�lHＨ��۴�����1�8�:�_iED s8F�� �6��ra�G���M��=���`;��\R�Mi�a�>!Nᷖ�0)�V�"��$���-"Ji	�0�Gp�_u��� e���]�?`����o�?4��Y�`r�vbcj�Z��\������UK���E�g�uqʟ��U�Ђ��M�z��l�I�������	�W*dr �j�o�`W4b�<��\��"~,�1��e�;�H���:�W�j*���n�f��~�T�}d�J"m�`xC}��w&�%,�������L(J�՝>�Cbn1�R����k,/��p�Z�KF�&�g๋����+>�9�� 4����8W�m�/�2�����������=+�c�K��]Bfm�d�GU�E16�I�ݼ[՝}{ΙZ�0#ĭVȂ��Zs@?�t�����R�4�z��X��]
���z���������K�B}��Vc�If��y��@�hgq�AW���H�G��j�v��FkNU1��a/!�������A�,�ί����F�ci�����ѷ����c����]�t��j��o���Z�Z���U����b������UOҞ!D1qt`z b_6v	��ܡ����ę`w0�勳�>��h� �4~Mڼ���@o<|��T^��1�*��#6&P�]"*��SK��|b�
^��Awa�(:1wXM�$q2�D�\�Y;�
Q\
�`qom_��ƈ_�Hz�꡹�)�)��,�7��E�y	ߩłׄ��F���0��g�˴I���٘��x�;n5�*�)f}J�X��8#�:��ԣ��B�EL��Zd�?6�O�,1�x���q6���ꝗ/3����E��>��L#�;��z�/n�1_������5���O�B���lgu�a�M>a㦆��`3�ݦm�ׇi���ꍆ�<��8S����7Y��!��'<<۽�V*{Ġ��'�E=�����F
ߚGl�-Y���mM��:�l�'�
<�Б�s��ٸ����|�(=#��!�3�Bc�W�(N�6�>��b%����S�0}�#�p�yd��#�c���j:���&�]?��
�M�q�Lo�A3�F2�ng��e�<r���mU�ը=O�K�2�Qa�p��) h����G����a�P]�o�t��P�h#
@+T���O$�b��~�c�`'Qb�u�v0$	Y����h�s����2�.����9O��N�m.��\���H]�V�,3G~~׎�i[,�(x�)�V��y���,p��+|�ҶX�[fC�t=�JH"h`����,���'��ݦLK��n�!�N��N��*m������/�DU���]���y��:$�9R=� B �w/�:�]�)�F�ok�o�:o���a���n�����0
�:ס9נ
�w��]����X���&�Z�G2>���vYx�_�&��Y��X�b���h�U���>�(}g�͍.j���#�գou"mg�`I�1�I�$8��7\���&�N���㑇��{O�_�uP����E~M����(��z���y����.����6vUCsM��z�=j�W@D�ڥ��	,h[H��(	ɹ\;�<�8�2�$�5���-���'���+�7��mӯ��Õ��rkAn�=c���<ay$����;\'��+B���!ғu�_�ԅ���ű۠�$IR�zJ��M0�z�5.������)i�LN����x�9��>Ga5��u
w#�M�o����Q�S{~9�N@l��O&忔�8��V�nu�;���V��l�R��|e��]�y���]%���δ��O[�gu���ⅿpr^'q�&�)dx@Y@�
��q�v�T @������L�(�#-	�9e'Q� +eO��ce�_��,b�l䒯t?����_�'-��|�5��x��o�O��⮽�7��E�Y.� �;�Jh�O�9�sxq�a�]���a�&7" ^���ϵ��j�4�Cְr#��qg���  ��nR�?�"6s��6�i�����KsY���f,�u��e9J�����&J�DQ��ڈ�k��Dj<\���=�(��0��el���ӌ���g�L�#"�$l�u��'��$�*ҁ��$1�q$I$p?_w�׃#��u[Ŷ�%�w�m���k�岵��d����p2��ZSA�C- ���-M��Fd=�k���˛ 4��s([B�پ� z���eSWH��`��>c/E�F3�5��Q��gKH����t��W^ډG=8�n��d��&��soXJ'���m�a��"��}n@6G��y:�Ogo��.�����q�&9���稘�F:ۘ5�{3����[��̉��uy�WMA������-b�X*�!��i��
"��
K����R�ը�ƳE��V��m�9b�:9�'��L4�*��*�kʒ܄:�m�V�~�M������<�����c���(�btYA�(�+���N�oFf&��hƎ��&('X+��4D������7��Z��=}�$��[��[p$��,�(F#)���D;�܂�s�i	��^�l;�J�~�D?'O;�=T��X��T�GtѼv�^xWj�#�]�t2���#���t��Ny����^�3��n��E��c&K�wM�̴�zwS�޿�µN�r�@~� ��F}W�ĉ�Q''y��T������U�#��mX ���՚��E$� �n����Q�������1Ӥ�ӡ��U��Y�$T��D��zM
��UZN��7����9��^L,ɺ�wS�
���4�ǴԄd��H��T;��)Ǝ	���Gb�l줦SW�r�NR]��%.��>�i�լ�v�׵�+��$�(��L�0w��ܬr3�o�]^�4$e��@�����x�`*eO��`.�	!�����%\4�/�~��b=P謸�b,
�'�����8;����Μ�#W�w�b��,�\G�ތā���#!����Um�Ky���x�0rf�my
�FI�׹d��1�:�T�*��(�{#�e��D�ȑ�N�Q���ލ�OC\�Dyx��հ/zU��)ڳMZ�6n�w��	��f�̸�E�,�ݣ�M7g*�"v7�4u�H3Վ���JI)1dbҭPX((��&[�lG���âF/���"���(&P�a:n�pg$��D4�7C�q�O�CB��4�t���Gߴ��� u�ɯ?sYc/H\��������O�M�p�ch�Ŷd��m]�YӉ�w64FT�m0L_=5T��:��[�}��#WN�?$�mO��ܯ��+�qB�1��h�["���T}����c;���1aPU��(6IW L��"�~�FhWIj��
�2Q��8h%�tMF���+���GO%j�<�=]$�Y��xr7�%>ԇs9c,�ގ�j�QY%�*
�y���d�Ŧ�����j���Ej���,�ۻ#	�sx�\X��w^�%G;{�<�&�5�NR�T؄>E(U$gR|"5B�]��B��9�dG�/@�(.L�Q�g���E�Y)��o����������%�ͱO���ڱ[4X��#�ڂ�wX�|�!It��r�f����eұ+�D��_{�4�˃{瀜#^1�|��?��0P�F����А��xY�d��xu�*\�*�ٖ@F]�����>hSY�Y��̼;�dJ��R����-��eLI��"�'�+�5s�|�A�p��Q�����_*���� �AXs�,��II��X,�}�`l��71�H��s%���{J�%��dOqAP��,j+׌�FS�KF.U-�� MQ�����N�9��o�*��|�&# �p��܏a��Wuw������xd����ZBS���\�e�b���zw�����g�F���6:�������׳���j�m�3X�]9[�~&�r	�m'��̬���:�+*]��SS�ިm ��Cg�Z]yi���`��6���u�柦�cm[h�&g��P�T�U��_	�� ���E��d�tk&z�����-�Z��"ftx�P(Il���H�;�AM���G�gv]g����C/R-�&����1r>�e��r7��1��t������]����O2C��Ȇϭ���~N�V=�8V�<��y���DR'_V����͉�?΁!U���E�B'g��ޖyv3=�����Fs��+t�a����DJ����޿�(Q����9��[M���S2ι$��m��g��M��[<!/�R�쩽�����ˁb��G�3�Z��9
-�|�s�I΅2���]n�|��ˍ�J�f��̌Ի-r�����(l9ܶ04�,�2�mmv��\edt&���ڂ��u��P�/���R���tq���=��Z WIe�J�!K6�m����riHn���Mc�ş-���E�縷�����zxȂ�8}%	#P5��b���{9�MFGBf;��D��4�)�I�>��b�޵��N�E�U\�Cч�g`�0\���E���A]>�kI�c���3��/M����~�(aɪ��ш�nm����+.F��wݠ��)��&��tH*r���7��o����3	B�m�щ������(����,�J�C�i�_���Er��Y����+�S�g����C��X�m	��T�|q�yn2��-����F�ʪ���QV�4-*e�sp�绫���m״���:��޲B%���-����ȟ�my>�]M����Zh�%bk��"�N�܂������w4��Se/�p���'Ӱ�G��0b`&I'm}������G�A"Э��֛{��^Iƾ��x�Xn�G��i����2Γ�p������L[����\.�i�l?�`���$P�`Q�%|?T}��Y%yq��@=��ԩ�ۊ�_ٵ��u�~4C�x���E �۸4�9x����Et��D�&?�0������]��s���}�����N�==9����tBY��I���S:�6o7�G� �L�"ψ���St�N�b�����y�r�G�26�!��<��o���exЅ�<7��r�.O)'�+c�*��/b*��bjTR��ϸ΂�9t���SVţ��V�X�U��q�>&\�k�J��N��X�L�:��Z�𤡥����q_i��Ӳ�Б@B%�>X>8+T����[�"[��[�N��_�&�>���3������[p�{��m��a6�i^�X%/W�(��A��( 4=�N|`0��&.kʺ�{e����{P���5�H�_^-Ϩ&��fq�A������E5�a,�p�S�(ǔ�T
K5�H��̐m(jU4:n��^���r8?��oL�Y~WU���9X8�g_�㠫�5��� <�
�h��qr9dO����[H�M�����3�]�Wg���L��vZ�B>bkP9:��2�s��Њ��P6Rh�WViw������64�Y��-��f����q�L�
	�?9GH�.ݦ�M��d�l���]��[r�x��Z��{s��3�P+��ݖ?�ҡSP�~4��Z�-2G�z
�H��?.��iz��l��u�_\U�su��ʝ������^V���p%�dr��7���G\�|�B2R��X(��e(RG u��-1�ER�f#>2#ȶ������.�J��]6�-�f�����j����;����9����u9��CM���TrL�P������ƄY�Ӏ,�
N�óLf�O��ۚ���M��Z�-	��d
�,��);�iQH�gJ�%?0^\\��ː�h��H���"����$o��{���}&��ŏ)��.��,A~f�Bv�o�F�_��������\��H���Å�V�E���������*��{��FCH�-��D��� yB�Շ,���%e�����f�R-�{7i�'��g8p��m$j`����Q[}�%%�i�s���=���g����&w}�i;b�@��"��!{G�4�f�lP�X���%���'�Mw�|�N�x0�$�w;���K���5K����y���j�m�ϝD\�Q���u���[���y��2���(��#�h�`xuj�`0)�X��y�V���X���<إ(������QM����b�[Ӏ�zA��!41�_I3���^�T�C�]��37/���δ餆ʷv��������xMQ��(;���S�٢�Ϝ�>]D�{��ʠ1'��o4�8kT��g�^r��nJ�	\���I�$>n�I�,���^���e�Eu� �����e�]Exn�L�bv��� j�;�:�}��h���#��izf%�ަ�/^�XdH���%���|J�m�OE�����B�ш?�������Bf7L�2�U0Ļ��҉Ö[��P��g �T�W�͑�n:`KH��~�\�9��٪������շ:f�W�@�{x�l1���k?B����,M!~o��C���Szo ��l���f��w_��`h�G��\w&� m��,*$@�5�<-�<DR�Ke8K//͕M̪K}�ݧ�팧x"k�)�"H\H�kr<B*�=2�䝫j_��E�d�Wb�^Z�l�`;$#��t��^ͻ�^&����Zr��쏓�5�����^���丼��� w�v����3����r1��:?��+�hd�
�LXU���=D0�_�!��F3����W�a�XhQSZl���ʤgE�% g���h�R޴1�3�'-��S8�ΩD��:�l�����5ɾ�x�����:����)�����՚�S?��f;��0�����a'��Qc�Ӓŀ��i������3�q!U�‎�9EO�RC���a�2�ԣ�'*vJ�p�2(�̔'��AJ:�xa�A�{��W�;���,2a����
Ln��5=�%S&U�y:�m��=Ο�@�6m�2����2�aݤ(-_<��F�Ɏ�}���X"nٷ����E�6�|!a��g��x��W�a��T�	��=A^��=١�oS�*{��#�oo�C����p�q9n�%z����Y�+ S�+�J�QcnJ:Gm�[^'��B"F�e(F� Nҍ�=��7�xѹd�/���!(ѣ<ok\���7g����s{�H���>�|�CCP��\��9}R�gU�^�g�גM�1���c�����ۼ�
�_Q���?��܋�|���K���d�!�~���D��ܗ���y|*��g=S�T#�=:�2�=����-Owv��;�Ѷ��T>�l�":*��*��K	�I�g�to� ���_\U���\���xe �S��ď�������f,�5��_���O�衠Z��a5�6[�w��%���� MS��m�8��A��"d�U�=8gM�Z$玭_D�a��p��4�|��54���*}.v��3P`3�&F�JɅ�r�r�L%�+�������p�	J�k���iq���YZ��f������pa�R� ��~��)�f�0x,W�^��^o��Uw;�1={� �%�D��WK��y}*��e����!`�;$ǮĻ�S�!�m�����|(��_�ˣ�&��K�f��w^���ˑ`��+}�v���J-�D�����B"�aE��^��j&~�t��#���+k�9�c#�[�E�5��޼�fj�3Z��oQ�0[ ʲ$-�P�Y!!�('y�����u���Ӻ"��BR��8�Q��5�5������M}�VuP���܃�i2��#vhCu�u���0��_�靋���l��<a���1F�}j\��ܣ��_1B9쭕�9��%6��@]|{<��Tq+��"�٥��9����o�VZ�������g~J�צƝ� j-��J @M�*m�9�Q����V����$�$=��U�>\��E�Ow��G�G|ڹR�Y��7�
� � v]rB5w�p�=�v�G��S4� �h�$%�ؐ���B�vJ�n��� R�^ћ8��;t�}m2�5Ғ�6\,�:宱������d5�3�-��/�L������I����T��N1���O�C�P����g�>��k0r���,���9�X��̺�x�]9�L���w�@m����,�jg�4��������:�e[� O�a���k3�'Ƣ銋���!��DH�W���8����ĩ�ׄA^J	�1/A.�_���|9�AF�J�OŷD5�$��`G�v��A9cym��٨�Q��o�G�2)sz��4��=��r�#X��4Y���Sx��0��3���ՙLSc�Y�"1����	s_`��E��'u�tzK&��zN�OPpj���a$���W5.Pc��@4gT��3��2s�7}\%ZHW��0t�T��ݜ u�P-���.���'�d���D-bT���c�살gϜ�X��ݒ�O������lz
�V��zىɱ;���\ﳗ���
I,�:m1�T��%�^M?C�W0�ϸ)�����V@+��"2��FL�6�
h�&ֵ�{�G<Dˇƫ�Mf���̥���yK�3�NJsgIT�4���T�}�U��Q�0]]s����Z��X�:;�s���Y�p��x���<-�;�k+ �xzX%���$ =�y����؊�L��^:����9���7����1!+���_Z�Ԍ�A��&3��2�w�ޔ��D3�=����C$�F����ô�B6��4�Y��Xc8�I�;��7�����O�- ��[d�Х��Y�!f�) s�4x>ĺ}vx�?�Q����p�o��'�ޱ*=C]۟�Z�A>�`$�����Oq§�.�2���Y�����w��;�9-�rS4�Y(U������!��/��Q/)wS�Y�Q�����IW�)݀Z��w@L����Ue��(��>�pg�'�Q�\��Z��a	iNW>Ep U}���:zW(.Uy�*V�[��@@ @���_F![��wR�&'ԲO���m[�\�*j�i��x=齃"�GP�h?"�7�5�t���8������/|u��/���j�w����
�}��D�9%@��4���F����fUK�,Ւ��ų읨���x��5nӸ�]d]�0����Y*��1��2FE?���5Mn�}�h��O���)��*��")�/^��bID�h�ԈPr�]m�zyT��76Bz�`���7-��%�yI)�bfԓa�j��,v�y�����A]�]ũFąu��*�#A�ǋ��*h��S���Gp�k�]\�T�%���w�����������I�	1x�e.0X�Q�Ck��*���+~$ｸc��pV�ƴ��"����=�T��k����
7�6�sf�yy�)~
�������2<���L�04�S�\F�p<z/�L�i_�kW{��LD|vS��/$���٨��bw�o�����T@�E�o��}8]�?���"φcɄD8O&j���,!PA�$_�;t�x.�OLz�(;Ns=���y��ր�]zx�e�����T^<�Y��j���d��7�xOo�~N�{��s,�ʗX%�/�F򆑎S��}_*jf����qA���*��'������7�_�V5��ܬ�P�G��]z,/Y�!��|;�� ��F�y�����U���kY��ok�e��f�M��]@�i������\�1�~;��:�`�lH<k����r�Q}�bM�� ���/q�U��?]P�OϹ-r+s��"�BGbmY����]1����oB�c�����k��/�:���%E�E������/åJ�'����C@l5;�4 ��e��^���if=0���,t����+Jj',�d�so�{Q�-$i������L:V}'M~���f#���$��A���]��l��O����.Ge�A?\�hO,��c���=�:��D/te1��]J�1�g��I+��Ox��� "��	6e���&R"\��u_qC�r��|��u��.7v`�S�2�O�ڶS7�?&η�6-�~� 8��b��pD�sLI\2�L�1p:0;�;�����jB-�)l�8��^
��F��z-(c9���_�/=C���Ӕ��|=��{u=��^I"�sq{�g�J�(*�h_tz/�_,β�R���a0��n�d�Q"��3>�n�W��7׷#��E��_[��H�]��(s+��6����&4���.�L��j�v�-�ǫ�sngQ^�ײ��׼j���BA#aHd`�0E�?j��lު6[��Υ��)����݇���NF���R��㶼^��,��1"T�*���+�ّ�h�‘C�����/s�M�
X��J���"�*�RJn��kڅ�.��w&�X:P� ���	�5�'/�>r[���
�>����L���U�}��l��n��J�w|�!�Χ���mC)��.)>tcl.�dio	�z�+"n��X.�ؓh��4��f9���:���Rד�sR��S;bO�����!�K���`%G�Qq�w�����K#���"�c��L���e~�W��?��gnb�Q(��ꀰHQ�T	�����<<̀a����`��^�k$|�4���q�g263t㔲�hH5����;�1E�R��t��lEۏ�w澭P������9��.$�ͻlɓ������#M4�h�@H�n���U�����i+R��^C�b�x獢��8u��u�픋pB��B��~�+ yYЉ%��Ԯ22�����0S2���\���e�R/&��:4@�"s�ِ,��Z�h#n���w��v��S�݃�����E��5V��6�3�
�ٍ&+�"��\��e�?����4��*J\,����$f��8��dduXj�fi�����os��{���h.��i�e7U,�.v�J8���@����^΋EɃW���.��t:	���J�ߘl�P?��n	�(kv(��*uR����M�0<�L��@�Dج�=:E����{�����M&T� )E��C�Yf���k��R�U�Ζv.��D��nG�k�u_�.U�m"�3���$^�ɶh/���?�uc�D��Y%�}�-I/������pXK}������[d6�q�I�]��Bk�v}��C���Q�∪$���-��J�f��`4���]tՋs\�J�$��dk�5��E!H����gj�w�}H��Ŧ�@Y7�x��� ��+Bpܖ,+H4���ʢ�z ��^ZF�y�ٰ������C*���0�d�@xҏ��+���(���ijU;T��JH���@�n�y���1�J��N�xO@,PB�?5�9J�����dW-�07�����J�^��Ɉ^T�K:霹��Jpn����h�	�%@�%���;IC�Pߪ�^���D� z1m�+X^����$	!+P�0�'��e�TЉ�r���UmS��)�0��_�uԷ�ذ��I�O�a��n�k�jOW�d�papJ���k�?�ѿ/�-䏇���;k\Y�<��8�8U�0 _�*���פּ�'ѣ�g���$�dۭ$����?�� ��dR�l�l�*\�l�t|m 1�SĐ�Ж�
ҌΧ���̡�fOp���߃k�r�`Y���˚�6�{���BQ!�e�a=�}�%�����l��g��[�L��@�"RM�����8纬�ǘ���˪��W��D�F��V^���%�1���6�C�}���Y�\#]�|��Aq��)ѐ1�"X[#0�0����`v���3�[]�l��ls�^�ᓺ��ӄH]���v����c�楠�o}��.�l�bfc0Isi.etwvHơy:�\0P1����;�a�du^�P3t.��}�#���?���Ifx�
8,s���V��:J��<�"�6���E�ow���{5�.Z(�sMpQ���;��{k4��
�e�K�`�]�筚ڼ*^�݋Yc�R��J���e����l��ȡ�E�j���|i��0(�<}o�-�9&r�{=X�Q���)w*�|S��p*�����;�ٗ+ਥ/|�G9u�t��VM3�8(��νB6oK���� U�=m
��S�!᧧�i@�ZZ����<�� ������������Hf���N۷fi/��Y�S�p�F����8�mI�hM]����N�&%2�aY�|�FJ���'����,�#��lŚ����ʴ�R����jJ8�>�gɽ7\
����"5�l�v:	OL�����L��!d�Z�2`�"����B�o&��z[~%'�^������t��}E��-�l�P��r�CpE6�i���SCT�Y���Tۄ-\���+�8���7�V�a��=�]�5(Ä�LuŻ���7��˵{�W����J+�V"�/�7N�P�~��{�v�E��.�~QWn�m�`m�$�=��n��=��1uΆ,g֕^�ntås)�E嶲��E.�`��|:[�1�D�3��-ou[{�갛e��*_��~��Q�h~ ��`x��iG
@�����-ex |�b2O'���N�e��-D��(��>6�QE;�v�_YXq�ܾ�(�_He����nui,��WaFhF<���kvlP�����N��]I�o��o���2�UI���Pʿ%(0Mq<��/mo�+5���=(�B��w���B䌻���{��7SՑ�|�ک#E=���O�m���T�K��x׸22��R]�����@�lx�l1�^���-�l©قZ�d�jD�6��kF$rI�e��9� �j�M����;�y����N*~˜R2�t���I��w;h�Ŭ�ך��ư��\���6�f3�H�
�G�\�lm�����m�b���h޸��Cx��f�z/Z��v�|Ù��fB�;�B�؋{jJLX� ���')�1���ն��2�!v�J�J��INa�kRz�VL�1Ly�#��!���������`�����1�Ӓ��R�W��J�m�LH���"v��$��V�A��D�Nk
�̡�_�_�6�G�mhn~'T[\�Fn�B���H�+Q�4"{���8��{�4&�A��}ZoC���AJ�F\�*��W	�,���
M�n�~}���R�{��P�D=GF-k9�Q��4T���dϲif��؝���B`�&Eqoe����G�d�<�4�Ĳ���~�tEc�)�V��|`LM�(�8TC���XZȳM3fsP��#�e����
T��Fj������EW���H��#�Y�tjl���اY�>�PM���7ӛ������<NJ�������+Fm+�/�c����H��h���t2����ڮ�1�\�� 
Y���2�DP��#kQ��G�@��Y#�V?h8JZ��;�vF��i��6ބ�զj�&i���[JCD ��e��3L���Cw��5��X�Ȑ��V?U^���Y����y���f#O��z���|�#"mG�xa7R�ɞ/�f�"�T�m�t���/�VN��8F�~żF5�~ѫ֪�zi�Qm�m�1��i�;�k!�NKGMlW��O�p�֡�̒P�~�ш��a�<��\�L����}����ɦ����Ҷ�p�P��ϐ!���=a1S��xc/�h�BF��x+�~z����-K� Z'٦�.�;!��;s�4t�D	ЙE�K$'^ɋ�I@V��� (-����e�%��'�s%t��3��8=Q���*�4��� ,�|FjI*�-��&1 o�8���,�!�ή6��y��M�8!��/�]��d�e�d�&�$��J�`����cu��O���u��?d ����}�X���2M	c���=IU�'��aW:���N�ਧ|n��#,G�������8}�ٳ�R �-J�6M�*Ȩ����Y$}g <f�զ��@�4��H����p=;35������q�K�<+���i�*0�(����|�|x�����$���|ާ�Ĉ��~,��Wd�J.X	�ϵ�WZ���e�"o��fM:�lƔU�����b��%����t�����.�r�����٣Ț��+u�~B�1AYv��Hw�i�<��i,PϨ��N�Y/ˊ�<�>Q&�NkuE�+��W�Z%�t ��E����8��6-��k*M"�9��L=|I�O�G�RgrB�LT���H�n;��y1B7B���(
��'p�c[Ku�u	�d�no�%T������UnUi4��/�JS�� ,]����щĥ�Y&���>~p��h#2+�����eVX�E�4r\k���~fBC|L���V�^���#b=ݡ�0����#%�Dq
���0���*�Q6�sh� ��椾�c
��;�	����rUw��J{VQa<d6��!�fx@y�y�#P/=|(Q䝒�k���
�?����c���N�s���n�H����;2{��.l�� ��X�!�������LZ.cK�.B�0�j����v:�iy��r�U��L�=�x�m�2Ѷot���`t`��G�� @-�%��$6�v�Zޠ{!%x� l�(^s�o��&��=C�\liEb��ܛ *1)2����d��3��(
��qX��(��z��%N?>_�_�N�5
G}�9a���K������������HG������_���y[_��i�%�����>�F���E�2o�������m�S����J�c+'���k�*)-s�)X���U�@x&��｟�b��i�������^�dz�2Q!L#��0���?�:-�xZ/���4�u-+h�=#ч"��N�=,��L�|Z�6�x]��p��)Á$����S����F�Ī��^�ϤOXʪ�)v���98�tӅ	�^oM������R��|�،ӛ�|0�S��`���ǃY�	/��"ky�@�`��9�<�G}�&��1A�����&C��qj��
uT�x��Q�f�is%��gs�������-�/'<��)
N |���i}R7���Ҧ�~[y��W,��{7	z�9{{&>��b<�9$�	��~=7��O�q}�x2Z�yYRz�4BnU	��'D0�����n�,ꌕR-�^M}���n��$�h�`u���<��h�?�\8Q��a��)���K�Kl�|���f~���zhh����ZlL��>��2��� ����a|vw�v�a*��	��˒\�d/$��!"���x�(��<Y���:�7c?�~��ߘ��a��]������W�7�|�o��3�W	��8��8���������`*��eGy��W����$����f5����#Ox���R���D�ܧ�V���}��	>&hq�˖,���J1q�As��1>S�p�@5�{�dx2� ��~���!�yx?O�a7�	�gѣ���L��Y�!�Ր>��N`h�H�\����g���T��D�-x_��"'��m�߆��O�0u�� 6�Ͽ�=,7���P��[��so�Ku.W�
�6� ]w�h�JZZ�Me�`G�2�O��}� ��t2zf�nH��}&���]|9%��i[^�"�I	ņ,�y�4��)��V
V(Z������wF���S���>�]��+q�H0Gۊz������}�q\��s��5���#�nf��Fx�����aڠ�(б�Wr^���=�-�Xu�7�	�L�m1��F����K�l�M+fԆi�>��-�R�0;b,�^���������;9SC�q0��{��N+v�q `>��[��\��җ��o�L�F��s^%Ւ�e���Qgy������G�6w܍,"ƹ�J3�|�d~s �@=Tf�k��Fä+R�w�O���z�>*�|tq{�i� '���V^kg�T��}a2�"��� ��<G�����~&�Vj��&R�Q0�Z�֞����D�r~��]�M?��"n��(�Xo@�_�m�Uv�I����W���t;���G�wNgm�>�:|���o���݅�[�E`�t>�9�,�	����,���\�	��/d<HT�oA�O?ו��Ɨ�p����=�xS�\|5:��ba.���ؿ�(GҒ�z�Bڕ)�̇O 1�ïT�^љhStd�ȅk�]3@�!g����?Ӯ��az��p/}p���Ex;�����vG��-L��4B��V�"�_G˿vr޲�+F���-O�c��G1Z�X�D8zZ����$���o(�C�\��9�x��$4X�TL�Ґ"�<�߷f�Y5�H�:�Ճ�҆$�&ϱLO�����#C�;�c�I��S�I�e[G�&�.�h0��*������42���gR��C��?.m
Ǣ�[0��6�y������~�ax�f[���=&�%,0�8�%͉��N�&��I��ȷ����54<�8��fg����_9K�"���a)�����1�|�ĴI�r������Gr�����:[e�*�ڭ�������㻔F)��|��t�������jVEgi�Ο,��a�������k[��d����:�}����Yy)�UM� �nƖ��3��+�9>���bd[�:�oI��%c�t˂c���0�iAaR{���nO<�����U�	�<�W�j d��?nQ΃UӦE���B��I����}�����N%�˽X�ۓ���������T3}�����"w���L���K�s^��U�����0�����5A9D����(Z� %����h���=�V?�3�k�]b��\l�q{�B�)O�4��x�'O�4�׏�Ų�P�z˹����Y�E���(�JO�0��8��k�'N��զ�ߐ(ބDv7zDO�V|BH������O�Y;�c�*�~���AEz��n7��[����3��%�Yw;��r�Z��`%RIK�`�P���yt�ľ�EA���^�����W;Hs1�zp~��
��S(�B�Z	���XĘ��^A�ac�g(hF�k<�:�ϟ���)a��zm�RA�s}�S2�2H�'z�09�������Ĥf�J�z#K�V�;�H`�g�V�)��_���hƨ��y����N����D��ௗTE@�&bȰr���T�s2��+�M��!��c,zZ���l�!{�R�OY�Uy(��U�]\U�'ʃ�'��
���%����~��%�f{g���
��n>�gX����`{by��ˀ�̐�RyNj_��h�E�"k�������I�Ď�љC�q����cr���y����:�*R���3��c/A�܈��Ix8��
c����=u��D���,�bo��eȭ(�����y�|Lx���T��S�����X��Uc� XfSɩ>�3�%�	���R��W�D�rX!P�'W�o��0��؜�]���U�.İ��q�T�̊� R�u��R��Y��	d<��_*q� ��u�x,"�����CU�}��Y�x�%��R9c��9�)F+����9~^f,O���#+r��v�V�tv�55x�>�Q�������p���n�m���W���u���S7�ĥ���E!͆-��U}���k��9���ha ꪖ';�J�Kx��,��,k�M}�0g��.�cw0���b� G�@�وs��$�����se�^�H�n��u����k�Jҡg���#T��0g[A��M���t�7�9d��ϕ�ًVdM�{y��(�O}tg�Б>d͇:�(�Eq��k8k�J��ճA[G�����(����ȫ]1`��^��3�k��3�~�0�ih���hN�u�����Ϧ Eyɥ����<�X:]��B-|&���q�ִ7�1�"���fR���J�
s|C'�<C�^�k�
6_u��y��5w���a�|ݣ� s��L�.��Ox1�2R����O���Fw��H͝
��-��7k��9��9�>����3/�����,�F��z	'5����#lH��ڕ�����?�>��4�KXc����'�^�υu�Yb��>�V�����r��<	��3j[�{)e:M���E`����&���<A|�B��2ɏ�/R���QT�;ӊ;_���P���8�XMė��	�?^��%��t�D�:� m[$�p`E�x�H�s��am�U�$��'MP*c���tZ0r���\u�C9Z!�Ҁ}��`*T�i9���M4����qe�Ѩ�܃a̔iU�c�Q9��+��u({�(ܙ:�mr9@�C(�4]�����������T�ٴ[�OL!n'uSn�9A���^��a��\��rv���l/O��u�Mh��
L��8�5����e.�e�ʻ���J��P;'e�F�kR�1J����3ܢ7X�$,�h�X,�D	�j4F��S�8��u&Q�/�E�},h#��(:.w���
{�g	�e��*�Ty�jlK�y�^
�(��"|&������Z!3��Ģ��So���B'�aMx�w'����eUl��9g���4~ ����g��9�8���9�'�V��Uo���s=����Ze�pYz��CqR�pU����.��İw������E4�j�e��>ŭ���ujb}��ζ�� ���?�a$�DFq�(6��.�M��\��KB��Lj�(��vS�(i�A�5.ڳ!R�� �?��M^_�����l�-��Ib������Y���=o���.�YLy���,�r�¨[�e�nߞ؆4 ȃ�}i��O蕏��K���NL*��Q��N���).*�ㆥ�i��̳ٛ[Ri�Г���e��J9~�.{\\�e~{ߺ�`�\��/~"�������XuP��d�[Q��j]&\�V��Y���n%�V+���E:j���+E���B+֜�6�7+" �E
�������=�m����8XŇ���[�?%w
G�H ��&�y͘��x���J�6�?������D��/��h���7F�V�����
²ȉ?��&Q�v��/�LI�]�]��#�K3�v��)>�g*��i�eMD-=��:qy��o��)�=�W�*W��D���>k�Q[�����^<&������O�p��r�4/K��|C�Ε����G�P���=Y���H��h��u�<E3]R��WT���$��H)y��"�+���߅gK�~�k_����7W��`�Pë�64LM�Cx൩aJX]�m��������]еx��T���v^�Te{��SD�`��y�l�ֻ�RHu��3ka��'z	����۟�^5�>9���X���������"�Nx&u,�F��ŚNi达�gD�(0r�v�m{0a���9B(t���P���ї��2Oq1ǌ�<��MC����y�����uC����\���G�>����v�ˤv�G�G�)~�M�U��Ȍ�b�	��f��o�d#�4��h������)g���ֽ���=T�.���[il��~��uW.���i�2�OyK����Mq)ď�<��J5?�{�Vkb�?v�2�I����H3#,��G��Ϫ�X8���Ix�	66s��oy%��~V	�%�4��zʘ��GC����jQ��6W�]��޺0f�0�r5V�3��JOz!T���_fO �V���)���Ύ��P[��?a<����Hj8H)�מ���y�:�"+%j+W�A6Nx"����*��4��(�|8���@�����y�w�[S�A��'s{��@�[���Q�e��DC���U�X#��co�N��a�1�*��9\Nh��X���P�� ������_bz�ͭ$��)���C��T�#�NhP�U�8u�#x��a���,N�/��+
y�̨��1��k��&�̯�E~)�q��N2|���L�WXl��D�c�h��X��
�+S���c@W��ʑd��Xe���!�.��^�E��]M�:q�pJ��ͫUjM���ի��#!l�B��3SO�0'g�)߈�;�9gY��-��� 6q��umm���~��T]��1[xIW���j~ت~�
�|���.Cl�� ��y[�Őc��1#H���/i��7TP�\�Oѣ�9C������󙧝A�p�?��ƛ]Y@~�,݅#aINtQ������{�ԃ���S;����VTp�W��w,��vC(�Tt�%�&�ژ�^qL�4��,����|��~�P��t��	��M�vy�Sq>�컞�K;�d�h���9�E�I������#�-�M��;=�p
���b��v��Z�sX�Ӝ0�~.��x$���)#������u�o�\ֵv�@����y���dV6-7�.�G}H 	p��(4��)a��/�A�G!�+����	v�G�q����T��U����RK� �Rk�C&�`�؎Ep،?�!F�45��'���K?}o�ft�s�O��j������2k�	�%��00�R����Z3�耾 ���S?4|�7�d�Hb�<d�-�sb�!��VQj|%O �n|P��h4�MB�aqɋsr��/RG}50RA�6����u�?/4���w��b8��{��J�8c�|PsX0o���[ZE��g��d<�� ��^z���K)�$o5z~q����a���Ο�t)߸r�y
�ee��?�ȝ�	��L,��	R8�a�d4��(�)�ᇌ����gB�����>W<x����U]g=X�W�4��`��J�Č-�����#�S]� ϯ�]',0Ps�^W<��w�Xk�n�F�Wk�!��R��&����iSE-�'�~f�Y�Lw��!���m��b!��e�m������B���BĪn�7�k,����;7�$ �����͈o�6S������E}����!�t�I�F�Klu�-HJ5�RK?�ޭ>��}M��\L"ؽ��Ca�c�=�$@~	�����G^(J^�_�ԙn��4+M�[�k�$`Y��9����HQ�Ӈ���BR�4�ŀ�h��kw���(�| �pN�1k���L��q�
H}A)��4����zw!�?��ٰ��υ�G���C�P@34UmqqS�'�{Ҵ7*x��朂*�VX\�}���Ed��l�V��<�OOD [��ӱ���}۹5$@�(E�MU#]���N	��w���I���m6�XhDb2��v��MY�r�B�7�l��f���"ɹ�w�z0iW;}qH.�!�>L&��~Xj���#��m<��"0+�:�P'g�S`��Ƙ�r��^��ӈ�}<'{�j4�'�L\���$bw�rLRR�c�p>uY������{��xi�}v� �x�� Va�(nH޾#Hh��(�WءRd�{�{e/c�g������M��$��n�OgJm�I@�+"m�)��?jf�d���b�t~9�_�ũŤ	���DV�1T�� ��N 3�nc4�D�����[���в���D�-.�b6�\�l	H�w����o���̶�E��9}m��ju��z�����R��|T�䱾�[;n��TMKl}���*pS,;���Y>8�����aӦ��k��zc��g�|�6�L�Tq<�ʀ��. �c�n�5���p� �Sć"��ݩ�z��n�,��̗{�Y�+�t�!+�F]�3z� 30-F>��q:L�׼�
�h��ҝk�'���j\��e�#���K-x^"�y������V��ۯ��E��,�J�e�䓽;�$��B�P֜��yP�w��B$�һb��U�<S.$�enZ�8 jOg��NB����&$LB��&�6~;�N��2�R�Ԇ���QȩꂽhSO��z�֗U��37�퍉��)T�FBp��P|(T�?\z��@%!yK�����wX�ڕ�}���ٙ�i?o�:�8�:�4صd�J�N��L���6T�;�$c��G��B&c�s��y/H���K#ژ�u���7M�S��+�Л�	i�����
����H�=%>��HT���y�^ч�kpJ]V���^��d�>�:&�}���H��ŧ{*�cB�7sN�Y�3�]�d�E2��
U�I�#�W�	�I5k���r�)u���R�(���{&k�F��z�x���i��\�j(���B��8��0m;a��v�m������/�6���;|(|a�"	ҲA���Z��+r��,ӝ����&�?_��g�G�G�	ΎiG����*����y�b-S�|��A���d�!zϵϨzE-��	���aj�P5��������/"A.��E��V��@��+I�9�1�7,1�OƔV�VҖZ�Md#(ј�������G[ʪ���.�g`�(��¼͏���	4;6�C?8��x�O @UW[�mc��W)���%^�=Bn��a�\�<5�T�	!}o i5��j��6��x[�!{����}��ˋl�oF6�g��������s��9�(�� ��������/�38��Hd��P�ҹ�-��fi�\$U~7R���9�Bs'y��|?ӑ�."ӂ����Ğ��}�*o�w�4�$������Ѻ�	t�_D+��|���t��r�J��ؖ}Ԅ��PGο�g��_�r�ˁ��cFL׷Sv6=��;�kĿ J���Ny�d�j׆��+@����B�l��kF�0(Nx�- �l9�%����.γ�ϔ,PU=���y#�C#�&�tŔ�h�/ m�4k_�\�``�C���h������>N�?��J�lj@��?d�0,v�tF5�A��O��[�Du\��r�Q�QA���w/t�+h�3v��� ����-^���C�}���=p��psƯ��c��C)�v�(s��Ί����#Put�w�=9��t7,%m$���/b�E�a�- �6�p0?�^�	�I��|pn��Uj��E��M`Ozy݄7��aE��RJ疈�J���	7]�Q	Np���@�/Mܨ\a�(5�y=�瀏���Pt@cgVW��Fkрֺ3��#N��m����v�,B^뻔��WI]G@����^@H�@���0$ɺ�zZjs��)!�8����#a�d���n��wZK�i�a�SkxqI{��x�R�@��BW�[����y2�m����i��R��b �o��
ݪ!�J�JĢ²�*�1/�MɺE�j۴+`���%N�κ�S �����<�W/8�-`��@-F�6��zP�����s���[Hl�w�'�~1��LX�5CE���,g����)�o�H14��*U5ȳ@��ZM?z�|�/�����YW�}<���kD�k@%��)
^x�LUE�Q������Cn�	�)"	�������d���T�K(���$��~|�$�����S;X��&m 7��G*�wP�dI~��m��D�#ו�)����ۗ�)`a�:J��ݏW����so�S	5�
�|]^�84�&�P�b�!�X~c���ع�YC����������D4XQ�%#�]G��|kⷔ'4�5U��T���s�	U�R�O�I��ﯟ������
�q����ӏ"��I@�:A�6��v�F�6�ִK�ƪ��YQx��=`(<"G���GeӋ�&�P�	�M��-@�~*�6X��MF��6�t���kii�=��gYy�L!���1�P��kf��ti1צ�ԡ���`�gm���p�S�5C��j�i+�:�;c���@�>���z<�k�9���\�n4dV6k,����sVB�&@���������SU"���"τ�4��+�H��
yж�����5oT���<hS�ѧ�9H�`�#|D���?ѬT�7vm"��dțA(�A�&0��q�_���'����#�������2��@C�U���w/'1����o�vۃ��XE]�+�_ f�脽JJ�D�j�G����=�D1����J"��<��q�P�`t˼���-�ݨ=�j��	�>\7�g���`1����������@@{�5�<��F�X��&+�W�d$(�u�[��j00�*󆹡�����Y�\"��x(|�Q^�٭ݬ�ƞ֦2h�yG��c!��NIЯ0�^_�r���@�M�"� �<�ݹf�ηcй˂�6�o� �I˲TB�H~���>�P1��6�sl{E+���`�ɮe��y� m�+z����t������(�&z��7wPw��uO����e�gU�Χz�c&��04�	��3�]TU�9w,�H<����򱴉?>s�ֲ�/�����cq�
Q�H�z����s�Z*�I�x�M8�	>��f|>�ڇ�n �8UHqd�%������]nF�]z��͇�!W>�lX�X��"zwT�2��J�Ww�b��d��谛_����YeA�����cl�֡Ĉ9� j#M�?���<�N�(�Y 5��b�G��bڍ"x���G�ᬅ���؃��1��r�+� Xk���%4IＤ���q�l
��L��N6ՎL��c%�>k�IW�Q�G��K�D��W,<V[�R�[����|ъ-�R�D����4p��Ey��91��yǀNo��L�c�L�U�bV�^M9r.X�8}�?à�nA�70^��X�;��3�ǘ�Ih��L�C��!��O�O��U�ԚɘXG~�DQ�H���SF����0I/ۆ,����X����
��Y�'$��eW�fT9Y���@*�����w��G�3��9�ȠW��Hˑ\ �zU-=��884h���}�����
�`�]�dw�.}���r"����A*V��ϕ��d2�����!�0�E`Y��|p�}K��j�+�����h��� �=��Y�LP�U�̖#���1IW�|�+?�1�1K�g	.E�g:�K��@�[T��o�«��3�u���L̄Bȋ�%W���o�]Q!h�����^в�c;���ψ|��X)��b篐�R�a��!��Z�)nw�Vv�=)�vV��ρ�f���9�*\}�Gٕ!�(^��/X�J�7������ڛ3�V��+�1貆�
3%�:�^9�t�~��@|�F�v����Slx �m\�g�It>'���ƉVY�Q��EXyOr��[.���]`���t"n�5�½@��@U�l�	��ƃ��e��W�~r�^�"w��0����G�b�?p[�-:J�>�{�MP�4-0N�z�̔!(͏�t��0�V��6���$ۓx��y�^��Whee.&Zf(�!��'����ϔ�Q��25XR�h�Rёuh�F2�»�y�Y���ؿ�E1��#qIYݗ��S��v&29/40({�˛��%�f듶9Ҟ�+.�X�ǭ��#h��ԟ��w�v���^a7T���,O�V�ߝ<&/71�Y��㻴k�f�<F�k�$C��B^��H��hZS�m�
�������=�Sb?8d:���_���-8�=��@�k��ʦZk	���_z�F7!����Ӫ����������8���Y�V���^�ﶏtxsѯ��� X�	^����Na(��%ˏ
o�p��X��k�JQ��1�e�9?X~����\��J�(;[�1���_=�L�$�^����<�s�p*�}&�B=��f�(j^�)�h�2
 ��#�c;2�$�&U+0�I@{������c�j�f�����8��(G��qe���L\Y��;v6��e��'\����&#@������u,��E-E?�j��12�F��MG]vE>[�Ģ���Ϩ��?�1}:�-ep����I\X��5EW���4!���nWL�v�{F����R�n6^Zi,4���	�{� � ��xa��@Tꅩ>��/pɊ �����x�� g�/��b��~��@��Ԁ|��/tC�\\�+��{+��ț^�F������އ�QE@&f���j�z̃�x�rslbO���Na����P�ʇ!��1��5�Q�+_yE�*7B�NïL�+#��z�%�7�F�#��R�*ں	Q^��[�PH�$r�I�d��Jc�nCݺd��u�ŗ��]e�����tvOf�~���Wm�3��M���U�������]���-%�ߒq�1h�/�&'I2D�"�d���A�2��)���INm����@#�i��((�:��R�R�_��(��1�iAEj&�(A������n�N�~�w
�~���D���;�DK6H��w�`
~�(� =L���UH��5?u���pMP���=)�+	k�m^�+Te*���T^
�sr�r+kp+Y@kU�G	�c��+��A��k�e��q$���"�!Xϖ�`/��4P����P��ա�mi�g���Ju�Z�>u�=̂�,=��yFaf��΢����C<K�O�s.���W6``�Y,��&�fnz)7�\�*yE�OG=�Z�W�
��.��;�Ó���(�_dK�U�Ih���n��7�'>��1�d���b?2�6��Bӛ�P��$K�~���L�;KhZ6���
��B�n�kPM"���*e�	4�,@���kMM���.�����S��y83ۼ�O�ǆ����ĥ~�=P	���J-n[�k;_{�h��[S��0&��	�@��U���b�*U;m���u~��"���;�@��I1�� oڙ4m�>min�۬���U]�D@}1��fᖬ��)!�18{O��i]ޣf�V���E.-}$�:��i+�/��ς����6��%OZH8�)s;�f�e��ȜU��y�R�����ܟ�Mv�4�k��3��DK�0��a[[1;�e����Y�F���^���HX��C?+��u�-B�(&��T�>�ְ�1b:!ڇ�b]�:?�ڼ�%Vf~�ȧ�u��M�	�[�$6��:)�C^ŪpZP�̀�@1O1J���P����
���9Z�f\D�*A2l��P���U5�\Pt���m��ۀ���JT�˼��P?@'Z�	$f�o�֔)�!S2�3_(���D͇M���(p SE�~�"�)R�d�݋�KMb�B	�N�"Ɩ@qpaa�ɡX;C�h����}t6�X�eVLV���&	r���F.�ž@��G���/C�S�ǔ�2C��X�.p�ʵ3D5Tȩ�ۏӝ��@�h�.Q�z㉈h�Lv���t���xE�&�m.D[q�楺�G�} UI�Ki�>\(����UM�g C�=��֢�f%�#O���j\����� �2��q5ӧ��s���Z���5��C+�óI��(�v+?��E8�����׍��8S^�/҉ZO��k���@�+@8��\:;����}iέhl��*\I��h�AzI�=����(���[f�M\Tf���̆��S:
�ٺ���0'�'��d�\�����k&I�C��ôi�\�bQ�ѧ���1��1���	��2����O	���CI��L�����0�c�j�`P���M� -�����JS�c�xc<�d��0����wO8�@��o�9�46�r�<`�M+����YuP�� J����� &<��0^�T!!B~�<�����	��%L��>#rK"C
U}E�}�[�`����w�ajP���gYȞS�B���W��������E��dp!���o��w���$�\�܂e��y��A~�9�:<���\���9x�J'��=Ӝ$FG��UĄ/�s���?z�Z���T�b�{ǌ�2�J��t:�<��E�N0rsn'�o�+Zo�X[��rx ��O�+�\\@?n�D����n�k1���b�v~\�l����С���B+P�*���k�F����_�-[fՕ��`�̘���7�����J8�t=�v�-+�%��C<��8���̕D��y��h�ˑ�v�}L\>�d`-R�"�05͊wHs�訢VX���@�y���֯\���nu�_�z����S�����������-���^��΋��ޘ*��0��J���6FG�
� �����dN��4GpH�#s�ƺwey�.�`��)��B�7x��*�rTM��HX`n=k�㧟�4�����-F8܍ c��4�¤\g���IY#3J}����pe�5�0s,t���/ 1�bʋj��>{u �>�볼�(��dļk<BMeX��Q)c����J�T����f�e�G��_}�<?ؕ�k���Ki�61�v�R�����MfӚPYDH�>�6o�߄'Sa�-qaḾc��t5�ƞ�`7��g)�Eg�7]W��_�����: ��h����r��6a���F�F�9�؛���R��qk������s���-0P����)5�N����gc���	3�R8l�����&j��[����Ma=��9m���u��N!�,�"Ջ �Z���H�_����s�֪����n06Yp�8�\{��8b��5]�����?{�����A��V��Z��]��tsQg�G1�CK ��3�3�pŽbǯā��z䩛"�ڋ���#a���5gQp-ĎK��]��Pt��������̹v�PI�$�<+�;���W�4옴���$B��h�����wQ|%y�O�(&��:�͋i��y�+I��</�y�S�yZY3m�I��eI�W� ���٨gF��h`���\�q�����m�dY.��y�_շE��08]9hT�{�p���0����i��s}�Vy����%$�@�Վ�r����v���3\�.�0�ϰSr��M��>X�a���Q��[�y8~���-���z��t�q�D��bj��`l�:�&Ӊ��7��P׽���4��W��/{��x�{�2y�Ɓ�8JFy�7��ҝ.O�|E���g���I,e���-:�,��_���̚A�bQ���Y�|H���@��ʸ�����ړb��G�ac��F��('�A��pm��$i{�?~�@�Mʓ�bӓ���C��ZIx�y���:���
ZRrʰ���2��ƛ�_v��	���-*�?W^����5~���6vx���e�a�=��-�)x���Co�ª�aZ�Bu@f�=GÀ��PE�i�F���p�-�.��w��E1C����Rp�J�T�]��!�TC`�kl�R��r���&0��ؕ@�=G��+�&��7��z�[�<bh�~����O��_�0�e���'/|v��R?��fߴ3g���������h�uݓ��,��n&��������#KY�ȶ=o`��WO��#`�<��P����z��\�
.���%����YJ�^��c�|o�o�bLI���N���֨G/�lq�QA~-� �isv��\{3���x�w����͊���pFW�H˦-��J��T���6���!q�!�}���i���b�v�s��˽���;�Z0}�}�N�}5���=���CLă��<���/��Z�8�!O�`���=��o�r���3���!S���-|�J_:L��k���p�(��21F�5� �L$��x�엹S������:s�}�q5{,F_pE޼ݯ @F[:���b������9�%�ǦGk�% �* T�3� �g�����C�X�`#�����"��d�6�]��=�+�R�*����ׇd�-
��Z}�������I���T��8�7�K{�acn�-]v��i`��V�cn^qKϭ:W�q��@��H�>�>%�����~0$w�L���&Υ�.m}�ԩQ��!���YN�!�)4�k�����
S���$i>��~�ġ@���d��%7�m~9���H��b��2:t�,��w91{��uD�uj�����6u�~7�GPHx��p�fM��oyxw�� �.�w��Rs�ppx&]�)hȹ���j5{�ñ���Z��"h<^� �QS]��D&P�XdD������h���ԃ�諢�vXRWO��7	8)�8OH��G���X'��V�~���5p��E�`QaY>���.���G�w��|��E���6b�q��ƙD���:��ү�1ᮀa�c/�A��l�.9Is��ղw��{���EP�ws�e1�?h�x�2/w����R+!�J�z��y>�:�"����=���G����Pt�`�WG���q=�<���R�<���x��ʶ3���7���[
�3k	s;(�5K�ƅ�)ס}8��S�{j� �I�ŊU+g�Ր�Ě�Ʊ*Z�d��I�Z�����^�d�&ڃh��萳��(Յ�c��;I����t桤!����%��z��u|y��vr�����%o~���l��s��{�>�X��E�BLt�e�%V�M>�Hcc�tE���W��/��߅�p�z���ݟ��P��\�p���������W[�ʫfN6�_߼`�rZDP���Y~E��"�ܤ
�lb;�p1%������A����2���s[�@���-[���H*x��c��>����64��ʪke�i�{ �_b�Е��(��tk������w�s�
D����������C��cQe7$������;nk���~>��F�/����8:]�ܴ�1�dA���<�f�֨�$��������|Q��H��h=l}=zc	��u���x_Eצ��H�ȕ����-/�H�RW��.�d1�e&Njv�,�(�^ ��|÷A�<u��֞��U�	��G;���:K���tJ�� ��hаU��c�N�8NT��^	ị�V�g�f����K��%	�I	��*�
ڪ�¬�Q=���̶e�ϼ��?��r�A�5��0�%�U�A��Cd4�E ��).��qa�j�a0]vZR=�f<������གྷ���̸�Mc#[��< ���k����5�F�w����ކ�ՠ/M���b9]���c��n�����y�)�7�xz�k�qJv�ůӘ�Be���XuR�i}4�LD8oC�PՏ�-���:�?���'_��`�{p��p�T�!�h���䗰3iȠ��i$�N�;�Ӣ�.�����Gsh��H�iwtAx�d�q�N	H����]B�b��<E�Jp�8?	���G�4A[�W��Ы	i�ٹ�����1��U��a�+6�v�1�Yz		�����^\��H��?f��.hy�}Ch�P�<T�t p���uR���Xu�\��t�����,f��G�#@��"��U�ﳎ;?ħH�I�,�Mݲ�vQj��Ҳ��A`x��P.���'_�&��GV�[�r��I�ci2�8j$"��q^J�s��z���֤�$��&����� �3~�|f��� K��eZt;{�g�kI��r���yg��6�&�^�v|s
��ܫF��	 �{�	���`>sɣh;ת۝K6d�L Xv�,���=���f&��Vҡ���	�Ac��1%9@π�����͖���5f��Z��|x�b��{��	�hr�6���� θ��c,l���o��-\Sz�ɚ5�ܣ�>ƣແ 874Bc��S�>����_�t�AAy^�uh�ϫ-�>���6.�ؚ�u~��^DA�[���U�0�v 3�(B
���#m�����᾽�M]�2_��dy�@�6��0�<� T�<֜SV���7�����狰�5m����mѫ����G9b�����eF|�7�P ��O�����\ng�uNn���z�r�'�.㦴��=�8��+?��%g93̀w��I��/�?�t���63�����S�񁭝n@�w]�_�`��������M��o�t3a
���l�=Zu�Ņ��^]&tG�eNO_At��EXD�%Gn�n��,jl<#qmRI��
���jZΞa9Ȃ��Rn���Ĩy^r6���PUz
¿���HO�;`��a$A�F"R���_�W"VD��U�`���rE]Sj��q�ڞCs:F�rI/E9(�CQO324n�mOު���� �g���e}���i�0�Έ2='��хrv��)/5��jU�e���P�	=#"͗b�1c�1{�ָ��j��+a
>���FG�%/��
�k��C
�YZ���-��5��f/^�U�;��2{���/�����L�Q � i"�	;�EU]�ƞ_��V��S�	R��\��)�r�|�uvg��!qʣO����]Ƥ�^����f H�8�LO�[F1	�@P+	B��z���, ]$�c�.İMs'�}�8�?%���f~s�-q��2��?������u3Je6�uD6�ʔ� ��������~��.�&)����Ǜw�j���:H�,�m�_Jd�'}5����������ْ���17U����ot��P%	_{�"D��\�I�h�R�;�82�ý�ù����h�E���v��m�'��F�Or����(v��9Atò��[x��N�8�N�s��H!�U��`�;a�Y�^�,�*��P_"����%F� ������(ĝ���>��F�h2χ[��UhG�.�_��P���$�*��38#~��94�7�B욿2�LZvq�?h�Q�*����뜨
�n��'.p�K��ātΖ�\>i �j�������- 8��u�X���!��pM@zrlǲ	Ü��}�����Rr_Z�B�r'p'�&w0�8Ⱥnsh�8�u��	�iu�a��,�׆K�����e�ܕ�*a��]{fWD���΀ ��c �7EDx�pq*��(�iލ��Z�g�1Uz5�6ƮK��d/��M*-b�4l�<�4E�͘AP�����#�����PЛXR�W�)��^h>�g���.������k��h2��܌�~ɓ	��w_nN�ƚ�V��|N�!�ړ\�?��(�ݒ �dm�K$�/iF�=9��?Rɪ�Us�z�*eϕ��D���Z�2�T���䣟�vՠ���(q_��,�8i��{���oD��U�����`*|�h�`�+�ȇ��V�x���b#�&H�X�L� �����!k�ձ��߼.;�K�l����ꆩ~�$uH�v��ϰw�1g�:b-�W[)&a��sۥ�/�E���n��D"<c��׺s�8��:P��͌/kL�|H |���&a����Nַ��ς����� V�=u����[�CV	�c�������H>��sj�j��U�\/�/S��Tɷ��T�3ǚ=S�������Q�s���HX�U�ZK��R���2"�c�q�2�Z,���^��s��7������i�e�@l���1�0z�){|F� \�����i�����IT�����7ٗe4[�q_(��Y
* _�rn��Q��^�2��^��^�}u���e�g�I�-�æ �Nz�*ڔm�g���߻n��$w�M�Q%�3l��!�g6�8	�s��m'�XZY6�Tn�q�#�(DQ�HG�]&Q�#��j���K��PC����u��h�W�]��=י��Y�u�xlr�3sNl�(��"��謢ha��w��|ɑ�]�>Ћ�Vqv3
u���
v�/�^g��@��弖vN1�Зp��n��d�+V��2����9�	�&8� @�;�J@���y��M��dV���4)�Zʁ~2�,j3����e ����]�VleF��GD�J�е���i�=f�:��+����P��n�J�"%+���K�R��Ke�F2U�G���NB��Р9Z�k�wi0x �"�	N�����'Z����Q�n��'S�d�v���zR��y��͞m{-�� �x�o���mb�eJa K!��5�'��τ��aUɛ=�E#(�wx\V��`D��6�w���DM�ݥ���)@�D���������
�'%��O}��Ҳ����sk�x�~��'���q�w��w�,��u,hx��Jm"��?�%'�@m��9U��6����f$�V01 �t?�P�_�w��ʹj��(R\G�7��([o��y�Aٞ�Y�e�4��/Q��3v��X=6�#�*m�;C�OT��BƳ����l�wkG��8�\;`� �����v*Ĝ>.�7�W�=�ì�m�hkL	�qr'z��=o�Q4,_��{4P��߷R�OŞ�l�^Q�����@]!Մl|�fpK��4PK_�M`��9�[�����U4�$����K=i.�kVc���br#C���6��@�tG��d���B��a��/���la}��{g�͍�\j�õ��՗ɑ�3G2�ű�7��ɺ��4�_����}'v`^�2�U\��
����ٷ��|�'�^�S�0m2��l��HM��Z�T�+��C���9}��p{8(S	>�yI�]����/����J+ްM���^Y�b�>N?���%3�^��d|[Ϟ�q�sX�X�c�٣�]�9�/���LYh-��~��h�JR ;"&��G����?�w�RJ0�Ų��u���3d;	�����:� ����#�Q̬��VD#�Q%ƒ��[@Fp�˨�]cL��g��p����� ��S��ú��.!���1$���>T���o�:F�"U��X,m,c�㡸{<��R*�5��ę/e�Ꜣ
L������_�����fՐ�@�J-L�3�><Q$��73�k%��A�n�1W\Iy�W�A��jS41�p�~iq����Ig�ך*+�(���Zj�ғR��NPX�9R%z��(�o�ڱ��m,Ob����;>�GD���5�x?Xa��Ǵ(Qx��&���^ӏ,�#�MP����YL��'�Z\n�}w�^�����'����#���F��[W*�^�aq,7�J������d�\M	���i<���TԱ�Xo���R�`�{c�rz�O>f�&�e�X8���Z��]awJ��@���ڢb ���״ie�3�j���哬�%�+rG� �~c�V.�͢�Iі�O:�A{?aeَ
�M5xʕ�3�R�j���2At:�b�\!52��t�!����hI�Q�	ɱ�����g;�mࠛ8a!1��nj5�����o���a=�N���3n�frT�߮G\��{e�aHbCJ?���c �����O:9���#���^a�U�<o�b���KQ�0����B��D(	_ALl�`"�0��?�B�$�H���t-�A���Zc�p�Y����\;N��b�!�r��U	C�02w�\�{����o�_Gotwg��M�̛�5�:$<x�RV��X�\�G����P���1�X����aNAt/(0�T�v��5�ԑ�1�߂eQ��㱥w��w �O���B	��S;<{pM�E�p[�s �E ��J��A�$��LB
��{�q���a|���x���mf)yA��2"����8��C{t�y�	J���~U�Z��&���3r���
Ŗt�&$�s��S�� �_/p�rI�>��X�")� &oN�T�"r�=$:\s�XU�	[J}b�Y#P�����>�e��Eh����zs9�am���5�zV{��-w�S{�����{�,mƅy�]�_�v��4���n�qj|�f���qn�*�C���d?j�4R�Y�D��zY�!Єe$�k
cQ�&{Ա
�'��|��T_\F�!�@⚂8Od��L�-��4A��	���Y#��fR'v3?/�*>�����KՑl؅3��Y\�a��^Q��N�BBrxL��\�YW�W��b
m�W��+�t�6m� C�u2�j��1l�L� �6~�aJ�N8p5L��p@L�}�}���C/��'�ւ�*��P�v��~_���p�Vޥ-u��� (�ݹ������T}?����m��2���T\�1��/�;���x A}7y���M{�0!K�w����Գ�[�@a����G��<9�e�+�&>�慢�+��8H�6E����t��,%1t���|\� ��D���?�X�����3�P��� �پ�~�m�¸���O3@`9�����:����b���,V�a� �(�]u���Ѵ8&�ef���ncC=�v^.'�z^a�#��~�nm��d0��v:Ax���t�FQ�/ �v�mu���}G�s� ��raG��$���^fLR8L��D�[AΧ�M[�&�OR��m5����t(�,�.'�w�t��?Q��js��!HIQ.��PAP���>tq�5� q��IB�֎�$@󱍧�;A;:�ʑ�SquG�Qa4L(B(R�L#?l�hռ�r��A�
�$�F���c��Rmz�3�Gq訫Z¤d��C���{�����X�?���S�m7~�?Ѳ2�7�#c��m���/M/ �x�zW�2k8��nI�^�$oX˝�<k�z��v��}�q{��U	��� �"�!��(doʋx?k*޻u� �	D��j�q�`�.LO��r�K�j�V�qEز=�p!݉y����嗪�
�jb%��E�\,N��y��(���l���}# {dt{�W��3o����l����?j��n�8�e�_�g�A-����ĵ�C�ms������k��Ҿ_T3��p5�Q�듟�樽��Q��p���g��x�\0}��Hw�)b�Wo�bG�ʝ5���e���1�j�4�U�=���\���;�n�Ɯh`�ç�P��S������55eG$m��ŭ>N�����4�ډ�Z�I1�t�/գ����S_]U�o۷qJ\%��ɶ��u0e�*y�ݩ�p�ꡰ�2��L��g��^�xW1����5���:ϭ�6�yC.x1N˭�\�JN����˪)�S�ҝ�I�ƨ}��J�HAZ�=�M���X�|y�]��,<N�K �B�@
MT'm^�zl�m%J��*%�a�O��vtQ�B���(�,�Z:k6o� ~,
a ��M� �(�9 O�K�(������a���o��
�:S�y��֋�v�l����9Y�cG��x���>�d��AX7'��'YP%t��u
�oA�{EI��-�@z���
���	�����~��!^ʜY�k@���E٧n����F}7ۥlI�ˤ�B���Y 
�����9�9i��T�{q�[��N���/��7~�G8�y{������!N�)K�)�8AF��2������Rf(�zq�h7`O�B4�C_��,��G%�y� .���W�s���+57Um�	!
��K�2��ݜ�t�R��h�"[�e���at��𺛳��b~	�Q���N��]z��~�.���j���ޒ���D?�ׅ��o����g��p!���l83���g !� �k���:f�������;���i���0zT����#Q>'�[P�Pҷ(�
&.G�H)����"��L\�s��-��{Z'�}���*��O�j;k�Hp�V�����9E���/�qi����A��A��@�!Y'"ӑ�b9+ X�qג9��p�6l (�|	Y�}β�X|���XlZ�^|�ҥ���������B����3߲\��#�K�����%��+9�5�����Ė"_1Jj�J;bG�;�Tʱ��Ihd�@
�!d�^�!K��S�����zx�]���l���ߗ�Ie����+�Ǌ�/;��s�a'p5sYZ_�6�Zc'f�8�pz���zޙ����^E�J��ջF�U�0��-l�΅(�<��1����t�ŷ�k�4Z;���Ŷ3e�*t��92�	�!���U7=f%�M{d:tozwjAM��!��;}��"�P`�i�G�!BU�K3��OL�^t�;$�Q�/Y1�����6��V��Y�����8󸼐�IAߵ�o����5�f���9��}�j��i2`����l	����5�\��i�-�*�Je�8������/@���ʟ�(ӧD
+Җ�=P�\k���RK�T�/c(ğ�N�7�h����j�y� ��0�>l�R§8��&���4R���ß��#��&9���B���_0R������'\����KUV��-y̶����
L�K�"X��Eձ����q��fs�3l�ڧ+��++��L�:�v��mV�s!F��J���g�:)�����G�u!㴥��|�#�*h�I��w��$c�|�'�өZ���t��p�a�kl���q��HQ�@��#%���f+\_���U���
J����i"7+���X�F�>�JR��ВZ���ZM��v��?��4�ѻ�sX�p���9�L
�l֔�.C��o5�@2���\��!�9_��B�V�SPc"SAH���i��6N�q��W�#P�K!��@����(^ʲ<Ã�s�޻\ȿYɛ=4<�7��#��·���,	���:uZxq?��"V�;=����6��� �yF8�K㵶@)�;��tC�YʶhDQ="��Q ���T��ͤ��I�mg� ��	E�:��0
Mya��m	(Q�� �������]*T# � ~-���9%x�������r�݄򩴾��(,�`2�b��@���ݡ�[��Q:�=]��*��Ԫa��� k<�UYo�N�`<�Њ��!�����_eN��.j�I=3�7�	�E4�#��Wy��� ��ĭ���,�,U�,>q��ZH�S�\���1��a]!
-V�)�^�,����e^+̟���|m������0?c5B�b�E��wp��ɾ�{���v�I�"��W[TO�P� 
����=v�A'H������J�D�M$��s�9�ݔTITUY���hno�([��pv�1��z�(:<�����(#�g�W�h\���0�������S�a�,.���ԡ�&�Zj�~�/�uL��* =��ɱ*W�*��]����1��Y�=-��WU����a��t���I���6���,��S��0}N=9c��уP\�5D� Jw`T�-> @�Xs��t�E��9@ς.%m�b����;'Wh���9aÔ0�Y
(��tn7�wQU
	;�/;�i���+:���O�tXu�[�W��<�f�a�OU���`T�e�`(L^[���d/XA���1ؽV���̱��̅���K=�GL��0�}Ф����	��j������͐\��0_(2�r% �+è>O^I-�����(G�ʌ�8�,������r��ם~1(�Ã�Q���E�A�-3y�����_>ۮ��Zqfǐb�gB�E`O�^01o��-CD3����.��8l�������n�_>�J2j"��JCX��݄������mNY�1 �G�K4��s!b��_�^d2�=ۮ����7���J5XB���5��
B�n�	�����?�$��Ju�"SR�d�dv�>c-VJ������l�x��DWR�QKuj"�������@kbh��"��w�!���Qn<�J!�,���%�4"tF�b33�+��N�ǩ���\:�.��78�ѿ�~��s�-3���\xN��DS�rD��輕�2�cA��f�`x]��<�����,�˟�u�K�q��k��Рg�Q��DRKaņ��:�[�|Wa8�QNq�P-�0�ͱˉC`�c�Ju�l�^��z�m2t��b2�n�C� �����A�w�ީu)��A��BvD��Lc�~�^=Z2 w�x8)7��ڥ�f�L��y�{�giuH	H���`��M	�E�m�>�x�ͧ��Bɉ� �����hu3?Sfl���ٿ�q��'�>z	����� oj�O�5�.��	�g��m��V��B	ZyF�U��z^�j����e�B� ���)�D	Q,�u�<����\�+�ƴ�F��n����9� ;?�n|��:SJ�<ۆ��uOx��@ϲ|{v�*6��n����X��RFQ���i��v�<H}���4���U�]�j�r�{2E~*�E,�%%�cد�x��Nt��랤�U��"�SȂQ�>�!`� q�0�x�$F��ՇB�Z���̷�[+D��7����x�j��H5���_rCd�%�� a�]5���^�[��7�,��`O�"�3�tft���+�����X�o벩�`�p�(���H��׺0��S��nK�,�Ѽ�״����9Yx���(/'-RĘ*|`C�6�L�Na�\�=��oq��Ǝ��[��c9ԩ�B&I���P�&S�τ��,^�3\�p����6���3���z����Q��KL��9�eS�,Fm;���Z���P��]c #`�q�	�N��ݫG��0,(����e�������]{ƥ� N_z�z:���BWӎ��C��dL�wg�\4hMgr�)U�@��3�\�g��4[�c���AZ�+��+ij�osz��7�|K��Y���)�}U9	�o�{�&�B�l�d����?uٖx������C�k�=R�%y�1~��݆�b��z� ��ը�T��1TX��g0\,��
���NR'�_��v��ԑ0Q�S������̠����巕]����N�>PG��줦� [���Z�����Zu�J�JY�bYb����3k�u�u+Y�S���9 U (RH�cG���w��������<W� f�E�|���)s�GȜ���X�6��щA9IM�2!��#���@ o��S���[+���҉�?1^M;i�Oh��4�[�)� ��u�#5��p���V����BF�q�����ru����[D�,P�&�����F��~˜o�ZKK<���R.�J\]8�������+�=���h�Ơfz�P�lKn���雾�V���,�J�'��=dD���0�5$����8�6��u{8
]xF>&$�ب��j���ozG,adv��E�9^�<�,�q>�N_�)�K{�yZ�ž	�5E�'%=���g^��"(�/��^%kAV����y������~G��0�����kV�2��YAi�F��o�QV}m>��<tT�ѧq��D�������tKG:��Ƙf���fQ�ڍ:���ڡ�����FU��S�T
���N�+�*��gBD��@�%�q�eF.�9|9��d%	]�	�@v���8���aN��dv�2٭(x�(��z�y�ZV�hk2�a3�81� �(+u�79F,�G��!�&��.��?�f�B~`D����y���b�EF	��=V�� ���Ʉs$�No�C�,㼪h����9P�Si��;���z�%5�Șf��Y�F�����Ã3<�3�]5-�}@}RQ�>�L'�:lF���e0#�H��W�����ɯ\��JW3-:�9l�'�O���1��N'ϻ��.�u�ּ�MO�J������e�hkp�.
�D/s�S>!)�Y�5ju.B��_'����D�qa�bS`u[,�C�<����Q�pS�UԒ��8o�K��K��[K̀���<�g`�!��7#��ѸSe���^i.{M8�wʔ� ��iWz�� ��d���S��y�}%���g��4B��f��S]:�f�wI�[��pI�ӹri|�i����5K�~'���Cv�b*L�!�r,�rJwM�I���:NB��a����|������x��N��!�c�/[2Z����|Lܮ���pS�Z|��ɑ���'�`
ylk����B����pٺ����Q|���'걕��i��JK��xs���]o{��l�ȀHP��*lb����@�X�y�?�'G������Ĳ��Í{��>\G޺C��b����yD�	�c<����x�����G\Pt��_��N�{D7��a���
�f��C5�̶�ļ���b@�D��cPE8L_6s�V�b,���Ͷ����=`� �ⴞ9���_�HL?L���5�����;�K�Uw_Ʒ���;�f�&+�?:7Є�&v�"���P�-K������R��B��T�:�
te;�����R���FI���Ξ��+p�|�ά?^��A����3�Rq�"'�G��8wL:�}�%R����;�,Ք��R�y��t+K�H���ZCb�7d�[�)(�"`�|�U5x�W�w��6�� ��\(	�f��64���&l���4�F~����7�{�(�l�~���%��:�C7�NG\�����0�L6�z4�O��6e�e�GDkz�sZ��eG,��Ox�܀��s@#�>f ��2) �{s�"\DA�9Y��*E׎/�>S����t�BMw�m�K~�)c�����3�'6rI�Wz�1rQU��(\~�-��딹V��bk���M��!��*����%��*�1��Ր�w�q�[����}�<��r3	�ǁ��������3'���v
�	�WTE6�&9�WU���S2��d�M�F����^ҋ�����n��§�&��&oy+J��o��"��䯺��;
k�[鳊)o��iVp����h�G2�Yݦ�5N�_o�dw���[7N�Oy��5��6�~�[�y��ˈ�,��a�wg��0۾V��* g!3�+*�V�u:dO�H �o*���:@u{͉>�cYʭCG0�g�d8�J\���GyDG� :|�CZ���Uy��L��ҍ�������=�p�g�]��U;ƹE���Dk�&Ư!�J[@q�tZ��Q�7G`wo��u�A�{��S���H�t�뱝[:&&�޹�ӗ%Z8K�i	�1]$��hP���8�>₉2�h���T�
�,���y���:����"�p"�߽/Ds]}�8�6+��s���$�9��q�:0���c�dW��S��7��{�2&���k�8Q����?b�ej�\f{��EG5ݝ���ǒ��{gn�Q�ښ��+��֍n5��(�����'ms��:�풿
y�$R��B1����2�g��]7ز�B�H���;�0\��$s�g���;���W����|$�����]A?d�x�`Cg�������3�S�b���{��j�j\�2o"ϝ�&�N�N�'����ѻ)e�F��`��dk-`��C^Pw���S����&���Ӧ|���07uu�g�|Γ�~��>ɟ�[��#/�+��B)��P�!��-r(>S#З�1V�726��JB\�P�0/'S��n�x�u��KF>_O(��p�)�N�ii�K=���HO"�ή6�G��y��Q��?�'��d#v5�6r�[�H�x��-�d\	�e�t4k��K��&H��f�~|��WbO$����^�f��z��>{���[�7c7�S�j�(�U�wƧ��$dYS�O�=75���r��D��'��������ʬg%L�(���uq%z�>}�L�F������r�3�2��O���s��.��ٶYj��d�\=��nJwa��r�?HW�ר�L�J4j�V�PE4||�?�_J��hw��m$E�.H��P�%#(�;R���Jgx�
y�U�ķ'�7��E��B�x�4�8`�yjgo�2^n�\3�	�w�x�y���L�N���g1��_+ �����$�* �$�1��ls�-�,�M����� ��e*�o����q���		��#����׎�Qk�X:���)�M��m[@��O��T��0�ϓ`�N�gj�%�>���ܞ�B��h�e��ł�{���)\P�B��`�f��}��a�$�� �X�#ֺ�}�O�t^%`�/��@"dn=�M� y��{���~�'�Z�-E�B�U��3�0!�������:!�ߏ���!z#I&8ұm����^e޺�m�hע|OF=Wf�-�����'2���0�g��9i?GD�$ݣ��<b���)	�=������pmhg�t�/$����|"@�h�}:c0�h�/���!�j3ˍX�ĳiPy%���u����#g�w��%�-��v�+��:	dO��C��$��4���J���l�-��I`� P��B�#
�H��`���D��F�2pʰ��lh��x���J0���|�C^�,�Ү���`Z��Pԇ?}�����Y~��0�Ƭ���K�9�]h�c�x�����qH�dȐ-m�^ĝwɂG6,-wJ���ԑ�Ώ�U*��a×1���1R!S����C�\�\���>'~i3V�����F���UDR��s��M�O&ӂkg�=j���A;S|��	s� D��5�ӈ</�Pp�Ƥ\�Օ���ՙdv����F�vH����z+�lGjǐ|J�Y�<�~��I����E���Y����9����֎���h�:|��~+ۙ��9R��IZ�f�ׄ=����Q3)���axg`r��kCf�uu/��B�<�p���@�|9[��n���/���"�#�F�)�&3xE��錇d�`B:�)3��Iϡ��hJ)�R<g4A$��ѫW̰s�/{��������a��� c�ׂ֙>���%��gvf����=��
צ:�t���A�]�/;~A��2Ds�z�Mh�$�Nj������)��EM'>)���+�7����kF{������	蕱d�'�d��')�3{)d�&佩?�l��pO3=j��$����V���h���*�1J�5�f�u.Ԛ3�g�H�X���'���>�l<�Ep�v�g��w��YR�q���3�
�G�(&m�{i%���\�
���-M]B�!|#�O�� �~�x߅嚫!��-�V	� ��r�R���|��dWeOi�C(�h���I<�e�����^7�1�r�7�m��)� �p�TR��f
��G\�u:�H�G�O,�~��4�O\�у��Ҹ�*@�P���ػH��-4w�ݹ^�n�(�g��r���O��樄�7��8��h�"���m�OMD���_u�,3h%����Bj
H�ǇJ�_b�lx������q����A�l�isd����\�I [�X�����`7�B;!�$_�Ne�dF��8c��3��&Z��b�T��� �$�6�v�u�R���*@,;0@%�.AFl,��d=�m�G�&���Z�lݠ�G��>֒�,Rs��0萫.
>t�D]�xE�e��q�Zx�M�s%De����p��	)�u��F�F���E��������9�T�$g�x]v�:��y9S/����YƀhT�DW�҂{s�ڢ40����䉕�0Y����b�#[��6t0�g��Ѕ������{�82retݯҫ���?H1�qMB=ʑڐ.�ٷr�8+m��(��.�N� �&:ڽ�/���Yz��3����)<]�
�g5X[KqDr�l��W� _R<v�C�{ă%3O�]Ou���/;��.��F�I��z�o>]�\/e����6�Mb�q7��4�*
��dG�aЫ�}��Snܟ�S�u����������i�!����>$-��O�-Y�~��tu�m�V���C2�ׄ� �P���G3M苸!���W�t�Aie�|SɆc�I�kb��4�/��\�k��c^����r4{��
�3�:]P������6���?J[}Y h���m{$��4ǘu:�B_���T��j����gL?KO�bd�K)��U�q�R��lf�k))Q``8ɕ��@�%��b���$�(�ŀ�����\�z����lɄM��v-��ŉw!��@�0/�2����<穠&Jw��0����r���	�>��Jg�����'�Q����\�68I���*�>��;X�s���̗%��z��YN�tP�╷�5Q�#�S)�iϧ����h li��nI�+����a�_��>�M�86c���5wdt����+�л&2�+3+"w@��}Cq��_�3�o�5"�ߋ_����o%w���lV\ �������c��b��'��d����� �2�Z���v��5z��ReV�e=��w74u�(h�\Y�fC�s8]��F���E<;�v0���4R�R���Ѓ��0F 	��Y�d[(�$ӗ��������G[��nr�<R(1���^�m$^����9��=f�{���e� ՚���*�^��t O���$�ZH�>��6�����zMF�&P���x�@�9"c�]�dM�pB�&��r�d�v�Ȏc| +���M���# ����@�uEݹ&w�*4���0����G�J�Xܜ��:P<�[�;%�h���k�\����<z\��}l�8OFO�ps�/�����E���t"{�8\�N��֢�1B�0+l���h��Lh�s�I�aq2Rd���]��BL�&�:���S{�uwG{�w��-�﬚`�S�Z����*����dd؋���u-�2%7��@��'�$�!��@,�WWf)�-�7-ՃB���M2�M��>��/ҮT�}��e�糿�>5q�b��M��8����~�o����h���8k�F��N��vkO%�G�+ {Fٵ��7��K��$0xH�CsgpG��~�Wz�'�{�Ji%Svy�d@���+���\��n�n�b���Q{��8z5�z���U��4께����0Q���f�,�,^"o>T4����K(���] ����6������1���i�uz����5���S�տA<u:u��K��L�B�1��C����
��ex.@�8p�t^��:U�b�c�hLF�m�8c��.��x��'F-�ÿ��LK�Lˎ��Bl "	{�^���gU��И��,=�^(_�������^��,����RWO*cɿ�������K�+�bD$S��f��x�4���b{0��S�����Cڈ�������7�Σ�\ö��:��Asm��[�;������Exg��.`��f �{���rD48�׫D._M����M1��gmW����N�#���~}�_�޹���@͊a�ȏY �Kor`@ժ�D��N�ﾩG�/Rs��D��$����A�a?�c$�)�mr�#�kv�d�~Ut"��h6�V��e�㉺O#6��s�'�q�A��7����2��@g��Zp�U�C��]IFn40iO�j�`�(��RI�5'@Dj:�tQ}�L�M�`��1(%2�����.%.����h��E񋜩����Wfw�d�i���s��n�i�*h�e�H���a�?���e�9�2�f{��Ec^4��UF�5ŮX�挨���,�������Y_i0�g�F���cB�'t)�-q���t�i{UG�u�خ����E ���EB1�Э��k�	������V^��儚��'Єv�XD)����
��aR��9��HCH�5m�m�
�d͇��v��wdv���r���9��@�
�������G��م��S,�E�1e?�\�/O��!CGy��V�M�����fO�����
G ba�~$��ć8����+�鷢1꾉�-���ݟ�A<^x;�`gt}�q��'D��>`�zvUM+2�E���Oqz Z��)t��1�ca���ݒ����>�Ճ�޸�[�H�1�9e��q�
=�1�"�aϞ%�*��mKr�\+=�R�Ł�N�`�H�q�]g{KYc��C���'j�����Ԛ�\�K�T6�E2c�g�a���Zڡ�Y��j������,�!�ar	���u�N*|�hEπ�P��b'��H�l�D^
�S��+KЊ���u'��uam-�V@F�S��3�&l_����_�L���
(��$�!O�l�)3�_;�S������s��<Ј��g=<�6�+d�cO
���R�)8�Z���M�ö.zSVPUN��!��{#Or�B�VhI��f0}�gpp�7��'Ƈ�g/�\�W�X���=f�^"'E]O�i�o��TCCӪ�,�����Y9�����x�<
ѕ����P�z9R�h��H�,[o/�ҵ�"�!7�6']U�7b$��c���C�b�����I>Ja�1j�M�|c�R��$�O�p�\{Cua1»im_����+��M�"�9
�t�/.R(�+��
/g��bh����v�O^�˦�in$���WW�>�0����N1������\)���2a$�K� )�$�tp�>�֑!/5w���a�6L��usD�2����(h`�[d�lvm�>e�(|���ҴS��^�����q�lM�I�H�D�a�$�
�K�Y9>Q�Ê�W��]<ݰZrU=;��<ǐ,����Bo����$ ��J�+����̈́�0_yy�뛣������%^`绹N9Y��Z�+VD��4#]d�л�l��j9����4�����*f�擠�HI�y6�9���`�L�>��,[��@�F/C�G7O'��5��p�b�]�>�Yd�jl�x�ꝝ��0��I�ʲW�hIP�FԽb �͞g	+|���������5*0�t�GY�ƃ=��[��>�0�A�2+���B�ed~���Wp���s�E��Ԟ|H$p2V���%h������,$�KZ�k�ޘ�*o��w�	�����;�J/�;?ŀL�7�E&8��@�yg�sWҺ��p�g���L"׊�$��C�E�7j?�6m�>/0�O�LOC;Ѥxjc Fwt��;̥
d��dB�4Z�o��ֿ�Y)�X��F8�\
�v��H�b�+��DI�*�#�i�qP"���Qz0��2�+Ŕ��޲���'M5t�J�Yʝ�x���}1xK1+�&�O ��䤷���.s%<Ea-��1�5�����P5�'�����"O}O�ӽ��Z�i:ɽ!,r�#��
v��!��ݴUप��4�7��P͒Zo���p�.�:z�.��G^�������⡁.�Y>�DPߺ���A�pS/��"d�n7�=���^���=d�
���h�5�S�x� Z	�Kk��u���L�'��Lt� &LQ(��7���s�m'�����P���y4tv
n��)�g�4~U��t6���Xi��;$S��=ߪ A	���/+��K��3�S�}жr(�!G�s��X��|�9!95��^����K���Wp\f��-�aCրJE��㳖��ZD�h�SA���<�E*�'.Mx�ꆁ��PXG��,bh��f�p��� ]�G����^A�/�
c3���.[K�k�"A �É��fR�0_ �l�~���D�;�YuV�1��bp1}b�4H� ԍ����vM��kz#\�Ŋ��]z:fZ�|6)�
b<̐&^�[4�u�X*׏�ݧ��-�M���4Ѻ���D��y�|��O�o,�`^(x�*	l�=��,�\~����VR9����i~=E�}���2�@�#k��v¼ܚ�)=`�Հj���=ʻ�"�H��\�K�9b��U˼i$|u*��)R���a�o[�R�5�0)��N��0ð�-�\i����VUT)O�JP���Si��/�>��j��y�^�niy^�����PM�����W�i׏��~�^��o4ƠӥGp2CO�1�¤5�ѻ�'�rA��>8�"&B�b�O^�)'bL�,h	��աP���y����I�����G�\ib欟��wU�m!!�H�6�D��Nm�=�7*T9�������@�AhƋ��(��_� �V�B=���l$�'���'��IaO��j`"����d��ݓ�1��=�_D"�X����-�r�<кX��8�<��~��+o!E�,U�J�9D�>���u�V�'�������{�I	�Av�L��꨷Z���_��X^��;���U*������NO͟��򒝁�@������d��Fn�@��>��fJ�^��z��6�أ�[U�A姘,�{�!�3�U!�EU��.n:ɣ]y�E#�a���`��ҩ��4���K��E���U�ЅH��g�@e΀Ak�H@�|��_�f��loe1_�\-�b���MXk�{nBrz�Z��-~Q�c�4�\͖�j�Yc��1J'������E�eA��$�k�8YMm|h^��Q(�6�/���6-�L���D�x�^S��b��"�_����/nsG�
�H���7OSss�{Jjް�r���p�Кpy]w�z�.��D�_���d�u�r2���&J������ �l�ko�,r��D�wծ���p@ܸ���عmdԳ�ۏ�{]b�@Ԃ�ycϼb��O@��#�N(3Ǭ�e悳��V}���ZAW0����T�r2ZE�-)�&�����ف�U@I����c,q~�K�>�[��	��p3�Tϼ0�(/��L� i��=�z\�~�A�H�k|�䲁O{�\��QMfX�zu��PG�ڈ}����P���,�����i0[G���1}Ϊ� i8OH�CܛN`p[�i�(���0�7:Es۶�ʍ+G��<�%��^�L	���P��nm@���}<i_g�f�xXr�i�rI�rt;���� ��C�|�H��� �������'oy�
9x2Wd\�њ�C8|�;���w���!�`잨B�V7̚�"��=��w>8��u�7\Of�.J�) d ����:|�g��J�#]l���RE�¯�.�e9�� �#�y���� O�>0���x@7YD8:o��N�2�h�E�1<E�p��w �����UmDMi��¢�dJb�v)
X���H7ok ���in�ڛ�E��$
��W(V�i�<
����U:��'�I[s���h�6 ap�ƅ��&&Z�J���9y����V���De��'̾Cr��2۸����聄�'!��WL�������-�C��>\¯r2 F��?a߆ʹ����N��W�R�հ���;mѡ�j0���ǭ�x�6J�N$���U�y�}	UBA�[b
�A�N��<>���wt�O��"��QG�\����@'�m�6�$�>��Z�]~D�E)|Y�I��JF~�j�ؿF���.R��a��C�(4�%j��9Q�Gv���g�b4� �M����\��jԽ�)(pO{���-K^è4O����6��2sn�S9 �۶��\bm�)9e>�xc���$�$��	`�T�U��,X���e��E�ad%Vq��JmQw`1&�I�q�>5�75j�8^���J�}ס뻲a/]�E�V	��Y�$�q����R^��e�~����&�/��R���o�@ ɗ(y��	�=��D�i�ug1ƀ����H�%�b �G��WM�-����ۤ+{WI���� d��+L��� (�P� R�o����X:��jFL�+?H���$��K�u�:��<**�%�Z�'�V����_C�ScP�cϗ�b�6��b�@��݂c:JϺ����97��k�݈�^r��hɗ]���s!S�>�P[�Y�=�� ��>��G[/k���ՙ���W�נ��|t��,T��K��D���`�rd�<��� =׆�eI���Y�d��rs7��5a�%����5�l�=֩��*�>�F��[�t�E-�� �ĺ������V�?��vL�4gxCk�A�m��FTe�k �,�0�}�aY�Y��HX� N~c� ��[�&��r���%ה�]�K6������c�ɳ�X>"z�#ҢQU[���>K�u}�1��RjB�w�J)�n]u���\N�v@�>��l<��c��]th�U2mIj�3(�~�������_�B���$��]9�(�ǝ�懦�A�P9łp��Yy3�J���4��Nyqz��/9��aC0����2I�]�hB�D�%�,E�n7w��~�!�>��ZW�F82ni��q����1����Zs����ٮqT�G�_��NT�V�,�Q]=%����mM{g/���p��bQ����ՅQ����K!����(m��F��ᓀX�'����y#>�MV�W�򮑓������<��J,*�F�W�X��MtԱ��E��X���莎ʊ��+���/�̡ԋ��:�YFiSR����J=|	P�+��1����I`�e��9S�W��~�恸�G[���9����@��!�bT�i(@�1j�CĦ�A��ї_�'���U�9�>�X� :k(��'c@y�:y
˟�FC�+XEF5bI
� ��7W��Wp�R�|�]M��r���5�7`��Y�o��;��Z�F�z��6KB1#z�����b>���*�Kgna{2I���b�T4�)��C�x6*X�,XY:ҩ��\��
ӽ
����`���,CcM�Y�|*+��mc��Ү���{3ӧY���<�m���Ij�ٙ�ڽ�{�ƃ���q�������ˌ��~W�P��ۑ�7"\�T�b�#[�F���m��j$�wor~Q�ց��^1^�\2R�1)^�02�S���T�T��r=8'���|<�'�0GT��� �����n��<��F��t�-�X�:�y� 2a��_)���Ps��#���p�Ww�L��b-��4ojv�E/��v�/GNL��F\Wo� ���(3������`�����T�Fk�W�*����E~1<y��l;��n5�֎7q��Ȑ�H�5�u�1��{\�*Ņ2](�,��y-�Z�n�'��P�~IR��	j��G�	:�����|qL�����o�'5v��
�� 3sL���K��c~�׋����㧴��<8(�w�����x����`�qqf�?�T���qj�."�n+	|�������Co96m�Y?d����@�R��J4�U��J��G�1H����Ovv=bV�p�-�'��~G#	d��A���Y���>,6�����44_�Q�o�o����=�ܛ�p-�
�5���?�4X�2��;c�z$�4㢜���3������3���Rqw/�o��-Һ���E�x(�ı��s�+��d��0�E���W��Z=�D�q^�z��}׭�����w�CBb"U>�B�w*�Q��{��Ӆ�|�[Ek��|�0*�=?��I���yD5�SD�A���z�g`��T�Y�^/�y�/p��+a���!hA!��K��6�Q�+�����TY�|OBqJA�ʺY���tB�u��$j�G��´�x�/R������z��M=kV�2����_K�����HS�)d��Fe���(Q�x���n��Q;��`.��j]�_�7߹��l���z��[��#@�!v�R�?�q�$$+�%|��%�ZP ԑ��F�ݟzS_P���q����F�-�����?�CI���y@�g�����t���vLQ�xb���I�ւ˭��Z��F��=՜�ڂ�Q��,=�!�˗ �O~��!�]Ŵj�۸e��Q1P�By���"���b�2oa3B��u}9��|� ��W��x�$>��>��/'�K�--*f���~�ʭ�J}R�!N^TS��p�P����h�����A�Qs�5>!��nu�sBFq�0-�+-Rm�����q�(n��W�h�h&��A5�U[�d�C�w�>hOf��f�Q"���%(����*ո��N�u��clGb�_���ǆ�c{ 7���f^��,r���f�Z+i%��b�5	���@l1���&P<�@x��a�븇;�ķ �ے�$��ޏ��؊#?�6�bq�{x����Xf��7R��Q0M##:��g֘�����WF��p�`D�tCڹV,6Oq������(ۂ,�<~]�	��`�oT�2<�0���hΚ�\Ķ��Mz'�V�ڡ����*�Q/PQ��Zz�K)���n�,�ͣ�P��l��bˆ8��1�GpI��/z�FS�8�2��z�������8 �:3)�4��f�&5�J%������v.�-�Œ^�|H��� 5��%Ă�eqҒ�߂'�ѫ�1�a�xZ��)���3Ѩ�pC��_jƠg b���[e��?��f+���tk7�T��0JF/��l�\D���G��5mzb��{�c����BÀ4j��G��x�v�Ô��^�����}�qZ�c�P�`{�]����{��l}?��!M�@����?\�'xQV9�_]C^C$m��U�PWp�%O#��$h���D��蓅��"�����D2cI���z���Y�����y���"�b=T�3������[ۓ7,�z[p��"�"��kaG�� $��ےm)�43t���j�4�5��/�؝0Z�m>oH�����W��ǳ犃'�����.�����X��Ha��l�'Bl��]���)����5t��E��O��U�(��3oO3���y����f��6b��|}��/�5"�.#ԙ���+��������%�/�5�.�{��{>	�tkV��r��b��5�-v&�N��� !F�y��M��Y��dD�d�}
"@��#��ݘo�z��i��?�
�����	�ʼ3�L9�}z�c\�ɤ�BR��U������+��T������"<?���@U��!>��b�nЀ�[C�*L��w��R�B<8�9��5/�G@Q�Z^^��d\�;��v�� ��:��^IvϖY�x����+7,�&�_��[LZ3�h,��֋�u���D�C��A���?V���4��5��1|��)�����qJ������Vm�2:��ǗB�z�?���=�]�w���=2����GwH�9<��q��U�+�!���vH�}�2�B>�0�mδ�i�mM�
q���|��𜛛c@�z'�~L��i�1�nߌ�;�L���>u4Դ��pTOE�x�9�����V3�-��s1�S�Q�F�*A_-�/�$�Pb�i�&���{3�T���$�b\�hLr~4�V��Oqc��mMN�"�G|L���TػH/�Սt�\�Y�kZI�[<�~`�ä�\;�CQ��E501G��r��:���q����G�����A�7�k$�Q
+�)��؊Q�N}:��!\��\�T����F��߿��ŖhjD���q�wù<������Q#)[����:�\_)�|M>�"Ao*Jy}���.��	��eL�<c��1���-.�r�;�[ȕj�u�|��b�@��X��c��v-���QOƧ�����7�� }-^O���5�K:G��+���]v��ۀW��W_��^�j�[Jn�[P��4���{��ge0����⋊�ء�-���
{�2sq�,���N�K��q���ܿ?/����ݓ}F�(���6uvP�I���F~�x�8����y���Xj/ъ���jГ�3P[�	ɨ�F��QN^]��b�fL&�� ��	�s�	��uM�}�y~%R%�Cʷ��k��ɧ�<��_�"�Pd3~Ln�����p�L�%���� h�c�	a|�(�g���]�2������x�O�˗@'����s/U8Y(��W�����w��۠WE���rG�\�L8�\:��凜����!�$��[����^��S�C-��+��ZH�o7����@ʣ|��/5�l&�����a���}a��Y��\
ѩ�4���D�}y�#�6��i��ED75�i?UB.���V�IXx�c�M��1��5U
�H����a�Nj�����:����z4 �GF)gV��
�.�7$�)�i��9":���.�y�S��S�����`���ȀCs%f�P�a�D�s��v%���h�P��|���'��l��a�Y���y;��E���ؙ�{�Bm�}���͏��\�h��ו畈vg�k�6����/_�r@8sd�l���;��}��ކ}IP��9:L�P�"�0~�f��6���?�r}R:�ٴ4�*����[�l�?�>H|����"u���k����!�rL-/	t|��!ò����F�,6"���M���ѧ�}@# 60���z��V��|�E���U^b4;7j� �!|�� 7i}be��j�Y��ukC?�Zm��������2�Z�}G����
 E�Ǹ���,-;���� ��Ĭ/������H� +�@��ė��9v��S�����{�C�)�T� e X�&s��6��UF�<�![�:���%j��C2�x�.$�&��V���U��97	�ep�aA�CaH�]�~�4�X��S^s�V��������RD�C�����N�����@		<�_���(��sm5����ɶ{���Œ��t"�K�x�=l�������%��d+a�}Q!�5$��d�_�r:�����P"��w&(�ʎ#m�-#���_`�h?�1�I��w.�"�"E/ۆ=N� :�U9�g�.y#�wj�޺5e�{�$�i��j-���� 0��K�~�ҟ�5K�B�j;>�P���\O���^n?��e%�c@%�A�On9B�x���%����O ��,�Pb�
n���Z̀%�A�b4M7GFF�4�T/Wa��0�W�F(Մ�Kv�ȼlG~�Eb�;YD��S�*����5��صd��9��
}�i����eqz _e5��"�O��
a#��L�K���o��I�D�d/(���9��"� F�O�5*V�>��f�nV32��M6�+���:R���%N�`7�E48j2
a�g�QeSg�*�2�y���4����؉l�*��[�Cn��2�F��j�����w�V=m���vo�ؖ��S��h�����fe�RϏ8�G#�r�Ͱ�)I=d��:@�d�X]Hג���cH&�w�/�Q��i� p���M)��ӷ~��x����Q�CV[֠Ϸ{Yz'��IGǵ����M�/@cт� ��^�����Y> ��~ƌ<o��]�
~���F��|��\[�%�RS�����j&4������ :����mI'��#Q;IS�&���g6c����/3�Q�<{p]��40E[6X��e���f���9�|��+�0G�@����.l��Kk�'��z`�WVP@�wg���-�� =Z�;V7�	���v���	�Ť���n��V*<�_���-�� !Qh$[�f����\�2�B��C
�.d*wS��ڦ/`S�
Q�
��f�y���\�j{y���bo���3�-���h�^\hސ��8z:&x�����y7���`�6Xn0��.�����se�O/Ţq!\�{�m+����kܪ+0잎� 2�F�a�p��;`F/��ڶ�P��"r#��q?T�3ˍ�-Rj�N�������i�
2\q��2x[�5��t�I�X��|�n�H�ߔ5��_�j&fح%��r���V��FoaE_����ԍ��<l.ђ����|et"3�<2�,�&��9� ��o��_������� ��E�U�?6*l�B��l�l�J�0�,Z�{��Q��ҍ���OW����Q����wyf|�M���k9�����qG��v��>9̢6�Sl8��VSvi *��M
[��;�E���+�~��S�!0�&���ɚ� �2��=���	W"�"ˡ0�ٟn����Eo���T9� ?�A�̷��K��Wx�d�uy������j�ރ^H���á^���dl�4��b��Rv�	�s��T�ew�j�)n }y�}�ٿI	�7�
�����jߩ�(z%�%jkB�qH��o���-D��{�Pze
�YUtL�|�T�1�k�^�x�Eop��Fw���]s�.K�(ݝ�'�dɭN�%	�s
F���v6���{I;X���Ö�dEa�������`mO}>Ϋ&�q��޶H�Xw��h_Q�M���G=�0uio��"a���[��V�J��T��uRؾ�����ϱH ��|_���SB	����\��Z%�i�'�ԫ��y *Y�;\���|!�8�:�Z���i]!��j+�}{��rC�e+J@�����o�oΫYcT!!�'뉂tg��z�$n�P^�@:�@*� ��;V.���3 ���i��: ն�uyiӈ�B:� ���!��� �M�T�hϝ�Wu��M��?b}p��ʵ�����<��3�n� ���P�n���M��2ip��>���񶯥Z�"���^2c�a���i�auJB�,oy���
�	UiŐ�9D�a
lխ�_�9�c����m�n��Ƀ��*Յ��_�{1-��A.���=��K����.y�CƠ����o S����<��lA�g�B]�����>�
	6�lK��{w9W9��*��l�l��Wu��%��B�P��Щa��-3��9�G�d-s��:�q.�#;|TY�`��+��6$rs,�+6��u�6����w����<�LEҴ�d� ��T�\��@�%Д�VN��Uɇ�?��}!� ЦA����k��\���:��e���n���J����[`R�X����T��/:/�	S���,V��k���P����b<?�\�)h��/����'jt�lc}\}<O�cC/o6��p��`�{,�{JN���pG����ݹE��FP�L��4B�ģ@�U3�~�nyXYJ���C�a1x�"����,�T�YA�L�;���*<L��n�2%��P��D�8���[�/f�(���ѳ��R����-�I~�d�=*a��l��ʦ�?�KL�k^w5��N���[���;z�&�@�7��<��aM1��69Q{��9���Yԫ��;$��	oT������PBh���
i	���k"P�:M���h�!鎷cz����{pԛN�SF�gV�i|�����+-�|��h1��q��	����kq'y��$���_�zUp��I��\��B$h#�e���H�d�딝:�)Ut�pQ�$����HE�O���JnNv7(~���=���,t��7�}�xu"@�{ox�B�����V`t�?[{s3>�T�fb�ٴ����c������O'���ľ+h�]m�ND`�[��U��R���z�0!������T�g�ͩL7 n׺��S�o\Q���$��C�14�V hhF�b�9k�3'�l�Q6�N��o�N�ob��J@�(�_]6@9���&IGLK���="�F�y0?��YQP��U�<.C7�oǇ��Ҟ<���q"�~��F���PH!;�=�=�8�㾤C�,̅��	�u�%�r�ͽ!-��w�As,[��O�PM7�U�u�����O!�	��f�ˍ�0�Y�A�v�T͑�4�y$�z/I�?7\*�� ���..�q�BCz��Y�(m��\�� �EF��Q8 폞(S�2��� �����A���~*ڡ��mك�=�9vf����p��6#��� ��Tqk�i�yf��vh!���t���4KB�J���o���������e7(0�h{Cإ���,��!��L)���p�Twõ~�J�"��AY���ªy����_�X�W�����5V31�t�nڐ�`e�^��:�4N ��Y�?B��ionV^;��)|ƥ-�̵�H��/�_��+������L O��+2�_Q�:��)J鉭�@`��;P$o�	��m�M�%� c�J(�</��z�F��Tޫ�_��Y�r���ޒ@F���.Vp^�||"�{I4����R���'2�^AMH�{c�_���h��%�no�dq��R,�$���g�n�#�`��V.�]^kC6Z�A�Tύx�J�˺Z�K!4��%n΍$S�����7{1t͞4��[�1R�l�vv�6s(��;�$�O�\V۴�E&��v��Z����f�����C �e�o)��D������[�?�!枡��q�yXU�)r�6�$NJ�.�+��RAڢlnsx��7I�q�d���3�)���/A_YJv{�)s�a	�"��<�dw{\Ґ�n��| C��#���\
-.>�O�w����N�_Θ}�dSB"|j p���Ē�]�S�i�|g$�r>2�=�X4�6�,#��[��=��
�x9FP�R�)�����u��囻�QĊ�H�����<�wRA�Y�H��Iw��	�]�ͼ�pFҚ'��eh��EdZt\���Ɯc���h�v�N�������Iy����Y��h �
�$6oq1v+G���௹��h]��of-z�T�6�e�b�P���͇+S�ÉXL5�\g�4�BR�q��%G�ӭ�$
�v N:���#C٨I->.��g��c��O�����<��V
`6J�7O�u��P�/��[hD�������xbqq��7Gԟ�q�#0]n�$�W�#h ��3h3=(�؜��௾4F"q\Q*x.�[�-��M�6CW�xV�+��=+ژf����1�E�ZDG��ɠ��(^���{B�A�¹��W`��5��@;ە�0�윺�K�)�H�H�hֻ�TU[ߒǈd�W�yw�-3n )���,|ݴ���M9_r�۶B	OX�+�}=S�=�:���$aJ#����y1O>YP��5��7?i�L�	!���©�w�(L>�]�󨱼�>�=`NF��{��!d0Ԥᢅ�U��r[�b��H�[�9�])�`��a�@���rc.�ET<��ia��+�!0	��ɚ/sL7�������ػ4�b�����A �����@�[��uU��d��g�)�
"0�V��r�̠�?���%F�T%���a�7��I�T�?&d��X���C��oSc>7�s�!����*-F�YE�$�T"�x!�f*nOY���C駲��	w��ze���H@�e� ���%F��H=�ɸ���/�\\��7����v�6}��x��h�,G�]�H�W� ��A��\Bq;_(�@g�2෵mV!�&[��7yS�tw8s�����q�2>B��W���D^V���(Bv�&���w�?�u5c�+�6+��S�b0�K���ۆ��>5�
�!�[����-%��~���n]���(̱��xYK�P!���N�~��	�V߮@����m:nh�0���u��d\S&6嶦�VJ��?��^��l`����d#2����ͻ�����B��+D"�M���s8(e�no4m�#	4��8���1���baAFm�ep�[��ɘ�]��\ss��,��|��=A�GK����/%�O�[�'mXf*ͭ5��g:��<�^⊴I)f︀�7?f�d�I�eQL�,`Y��&7���2��h�f�O��� ��J耊��M�m��H��M��f�Jv�i8����k��n�������~�5D����P�i�D�0��3@=�'mg*e]�8,&Q�N���4�����k��b��r^���Ѳ f�Q�m�[��vF�d�ىU�JE��qb�e7���� F� ��$�7�'�-fͨ��t%��%s�����}&�O4���M�>��0%2=~�oN�Oy3|^?!ؕ �f�����N�0��:ƢG�00#�+�D�6@0�?٠y�s���0��s��p��[��F8A� ��"
k�7'���4J�N���u���;�f��nUz%��۾�����l(�M���9����>1٭r=-�N�k���_������Iݕ#�N$����OCT^�J��nD�����~��Q����`�r�� <��dCҪMzrt�P�6!��(8��~�syw��cg���z��J�$���"oS����}�����:%�p�iZ�ڊ(�&�������SXx�[<�_��~>7��p�X	�c�p� Е�gn"8�oP+�m7Ta����I0n�?�YZ}��̟ևK��IK/ʖ����� �j���a6�����C�ӻ+�B��4ҧ3�;�DZ�(}�<\$���d���&�)1c�����ˡ�p/T�c�^G$�UV�%��(�[�nA���S#�r�P�顭M�Q�v��[2�'�k�o!�n;զ2�mE�nɹ]��6��@?N�gQ@�f�/�m�V�|��!��/���PM�#j*P^[�J��/�u�k�q�% 4�7"%�����I� �c�EDK���U�4���.���pF����@�-��~@dVԯɱ����J�F�͕ �O="j�u����� ���gA�$��6c>uu����2��bͧ���)��5�>D	@t��[�gX]sR��B�j�+�J�ڈ���gELԫ[�6O6jp�%X�O^<p����>�I�<�Cd��{c���١�S�T����N��)�X�栥�y}��wyV"�?�3-;��fc��� �K�f^b{�I�o����������D�c
l�+��?����D�q@�ay+��L���sx'��d0oeC�	�}���\|�t�t����7�D���rv'��Me�pՔ�5 .��C�c�����w�Pc-Q�������ڍ!ƺ�44�V�bt���C�D���^�N��Ǵ�XF���*��)���=u���-���Vr����N��P�A�=�xW+5�ܔJ!�o��8�?����m�V���&5����i�5ΙӿP��1֮����$��c+�JT"�<ʶ�"��&Lzz��s����-u�)����A�7s7�|î�](ED���Հ|�m>�N���,�@�$�@�kP��hg���I��Ӟ�g���hY��u��c����(7���)&{�>+�y4�����^��x�iSZm��"���o���b�%y��O���-l�;~7�d-�����f8����O�?�� qab�hs:_��&P�OѾ�ێ^]4eA�/;����z�/�3�%�M%��dk���UERؔ��*su�N�3�]�'gf*1�����,>�x����oɤ�h���1�O���0���1��eD�X�f�%ø�až`<��󥂌������7CJ1"ួ�M�L���m��?\�A3�zf,��V�����á�3ĝ�Fv89��|z��%���*�AkG�}<Gm�~�;s&$��ly.�D#�c��d��r�,9��2w�m���1uՉ�MHf>B�\7<�F��3�}�9I�LPƎ��Jt
21�J�����Jڝ�הmU<+��K�j�$l ���6TT](��%�m5�;B���_���T,�x��*�_!�0(�
�WB��??n>L;K�ƌ�'  _O��}�U3I����SCT���A�2��G��ȧ?Թ6op�Z�h�qs��M���r�'�O�9�.�|U�&���Wk�Uf�/��ü�]����J7��H@:ZC�� .���h�$ʈ����Rb��p>��V&�\���P�*�K�D����;��xCT��'������{��;����_5Z_�y��u��]9��#QA��k�����)��xӱW�B%���r�(}󰍗�m��4Q�h ����8A��r�b���l��=g�zO��)V��Qqs����s��!���W�]#dR�wQb���Q�[��� NzCG�2���XX����v��Q��
�Xt8����4�C�?�ҡ�����������ё�8��U
O�ۅF*��<��H��*h%.�#���5N+�sX|�g��u��튷+u�λ��ݡwK�'Cg,A�/t�TNS;X����.H�B*�EU]�����A�a���
!�Yq��꜍.R�7f�I��-��>A��㤡�˚U)��4y �(��=�+Ƽ?����o�h�d���;t}+�C��`>�ؘ�
s{��ܪ�U�yA��ֿ5F��^:"5�n������(g�}�>h�Qn�}���LW9����#TF�����O3G��~���<��:�+<��U�喝 ��|���bnڋv�z[���ΜD	��:��{b��b�#��V@��)��q�/LDn�}&n�P�}4�+�Wt��`�`JX���t�&�3��1�m.�hXB���f�G��V���`�q_%�Pr�'|�v�Y�����IEz>��B�D;K!���ʊ:{�A͕�_�����$��B�g��0�Nw��A^���:-���p�W�0��%�&f���~�oQ.�'7?��^�f�q$�#���ؐ����G�Jntd��l9�#J=�f.E`�pMB��	�Q9c3�T^�W�z�ҧ�yF���˶Ī>�	𥴎,-ǿ<�AV�q�E�ʼ�����J�)w�t�5��2ԝ�C9	�UV���s��x�,�{8��V^��	�^aB<�wm�雞n��{��䛫-�`!y=�����Bi�J� �f� �w:�l�LQk>��(��bD�nC��T"����gG�a:�A_,��(q�u�c���1�ȇm=|��Y�n�MWѢ$V��8�e�hݖ	ꔏ�h� $���I΁%�����K_�b��{��wR"PS��r�#&.leh�s�.�f��Jw)f>�����\���e�-K�Ø'a��ڕ���X*	P��sq�L�1�>T�l+��ۄ�*�kv��b@��<��|덎�."�2�m�_�U%��
")��O~v<�<憾Q�WN ��kg�dp�Md��.,_�'Sr�QLi��
��٣yN�S]�IWu���Foa�e�"CF�(�1���G�~�ͳ�I�@������8k�r��QÔ�xA�	�5���,��5l�sA:��pS`V�̦�W����ml�L���2����^Ki�A�XLz�Uj��b�R��j��V��ֶmV՘�zvrfhh���m�P���&5
���1t �C�[b��'7Z�O� ��p%Ra"ş�8�/��q�&���ƙz�X`
j�>��}�Q��ֽ�P�Xz�[8*�BC!�J,.j�p�W�7�U�`��p���:{��!)pzc���˹Q��V�FkPy��P�M IO��Nx t�i2D3��F�;��%h���z���'�S�ҏ}d�����6���	f�d��U��i��+���حD�Z��E�[+�[{/���!^���R�����aΩNEϙ;��J���Hs�o��&��o�a���i�ꎏP�MŔ����¼bD;g]����a�
�+E`����v��KT�ˤ��ON{	u�[�K@]���_dnЬO�‥��|y�g��`l)�8�=כ�[eI�����
�aT�vC�)n 	��s|!�=�4`�`���3���q�����BOt�ê7D�-�C���JFGU�u�1=��s�޷��9Q�P�"�?r�v^�en�������7
(���{����L����h���hh���Ԃ����ԝ�$@��F���+Y4�z�m���~��v=fX�⇯W��m�Js5�X�u��륗E�pθn�k��L&�3���kP|�Ǎ��v�Ս/�>3��Nl�h�z�N=��#T��K�#A�lN������e)��ٗؾzm����e�ټ���Hj2GZmJ����:������W/3�����+�9e�����X1w�|��t�)@p�����_��OX��Q�E�����͔��5#�.�t����KB?K��ը� ����l� �ɸ��;�MY��*�!���s���_��U�I�#;u~�#d��_��r��+�W���������ph���~� 44&h�Bg�݊
�2���/�����j޾烁�/���弧R��!d�s��'�l��������ٍ��d%]�0����l픸A���E`Ø�g��iTmRF��Ř����� ��4����߻��-:�|̯9���OT}�7�,Y~Ɏ���d�������
/i�9WA��e�X��
���C��ⳁL���]�?W�"������h�|{��e�r��C2���3#�3�eX�$�B([ fO):�m���q�V���Yp�������J���t$?�?d(O�2��f�J�y(���E�:Pp�4*_�@'	ƟR�8Ԕ�v_ �Z��%ݙ�pY,d@Qj�ǜ���"�Zӱr�@˯h��4 S�@ЦW�qڬ�j�7���4�n��a�f�S^4C]���fB��F�h3,,r�3H���o�~.�Z]��C�;�<�%WI�/��� �\���$�Vf���mdJ.���!�ق�/�\'��Z(��L����,��q[��e�.S��8
�v�������|$8�d�.��yF�����fK������B� ��dOP՞鋫����z���3͚mo�$��Ϻ찲l+7Ȳ܌Nk���i:��^KY��H���g�?F�U�Ԕ�pBt���e�u��C��Q�-�\��Ȓ���/�
͕�I��N�`2�{��d��n����f��2�Wb5H.��~yY�o�5��qu��!��@Z�P���&��i���S�������pO����T�ԫ��+�]�o��Pc�d�b^T�"�U�	���{�W�P/G���P^�q����2��;�U��]JG�|�F�8/����Ƚװ<'?��.?��o�<�Aܭn�c։o𤋮k�����6�v��� �L�ݲR'�,c_���0W����X���0a(ݴ��BLP���9ڰ0�i�]_�.�@'r��x���[OLL)����=�f'HU{Q�0)���)�d�u���"7N���G���'��'���/W^��8�D��_n�M%���:LQ��
aB��چ�풎�:�C�/lew1Ve�P{kd�#���v~>���@+�B$ꦏd��~*V�E%+ �!��
��2>�����bw׊���!���
F�M�����܆���G��l1w4�O��L�[C:;4}�ب8?l���~���K0����%_6������Η_�扑�A<���kHn<�ڐl�U�q�&���Z˺=�4��r�\g,�jʹIFK����Qc�x�o���;���j�1Ǡx^b�˜�����Lǅ2�2=����̸-
&����6Sr��)��ޥ�m�[O�C-�`F;qvLt���i��|s{qD.�i���B`�cH�+(�cR�L<�����S����.�Q:Rg益X*� ��?;�`�I���/����k�d��<���t�0�Upg7Ddnช��F���in���E��0@�@�UP���%O�އt4��F����❓�Xܭ�:Y~ըdZ�}`$Y�[�Uo��n��bcCϢ<�&r<�N��5ۚeM��-~
O�Y�'�Bx��{���!�O�2>��~�w�u)r�%���Xd*3����iL��x��$H���R#�\B͓f����>�Cp�����ҫ
���dv�&�[���F���^d�������W,���=_%G1��ۮ�E��:�����9�^9��m�IE57%�?#Dd�0�[W��ݘ��&	.gx=
\A((a��TU
d�W��ŴnP��X�d����=��6������)f�+�r��|�^� ������
T�Җ���m�M���>������B���pk,�Ϩ��g!�,����5s��&�QJ�-%���97u��Π(#��W��(5o�k� �}���I�����d}5o�Ŏ�Zt)	}�y'��^���V=A�
��|�o�ueI��JF-{ۧ���������I�?���ldzn�
O����_l~eZ޶Iq^^&���BkH5 O\aĵtNl�
���u����o���M���t�qإI��;^y�<��M���L�����MA��^w�s�3(D��W1��[�]��O�Փ����@2K�S�>q������u�jx�*�m14[�B>.��'��m�#&��B%�����¯@|G���#@Q�;BG~x�e���}�G�U���SŌּ��}��	wz�
�¶�!F���y&/)��_JnHf��Ϣ�d�3�<���UR�5�'L��g6���}����>�q�j��B��T+�u��b�6PS�ǩ:F�������(*��M�w:��/BG;��e���Ig(��qҙ�-����2 ?�܉�r��Z5ڙ'����=�)�_�ȷQ ����s�%�0��)'V�V��Lp��ȈRQ�� ���0�z>8 �U6\q��n�UjR/?��$(��#�U����Y-*����`�X� �B:�spç\2=Ku��}D�$�5_Q��a�*<��!�s3�b��,۩��P�ON�A�yɢM���堭�j�;@��`�:Բ�'�J������T���{b�A~���	e{�/��,5�Q�R�<q$�yc���%���9��r��b���������E+cO�,:`hi��yЃ]�5��������=�)�C�Û�T��VpA\gQ��~N4d��,g��]6D{�kq�נ���^3qU�5��@����q��}׻\�U-�7s�zx� �b�*bpd�j���Mk�@h��� �1Ú���P]d�27�J���J]	H�L� ���4�V6�Ir<���I#*�jPj������j����1_[\��������㑗�-Ġj�8��m*�!�F�PJ�k�/����s�^I�i���v@�$8�~h0���@�n�%���T7 v���_���p�zr�x~����*Q"�#�oS���@��|�"�X#�1W`�)�1@�W�CR�9�;뫗mr��Lg��'�뤳x�t8���V�OS>���^i���Pu4��(�SG,�I�O^�I+��B�#�~�F�3FQɯeh��/�}��d��f�o�<�*���-;���)��p�����u	��_�"��Ŵ�Q�0��;D0�Ъ"���|%l1�o�6�P!��S$�[%�<��A��b�e��j��߬	����`��Ei��h�^� ��a���P�W$�!/��ƙ��[.�����\A��5o���Jf0E�
l�r�/�6S�4�0i7݉CsF�g���z�ݿ,<9�6ir�4}�6������h��F�v��qM	.��*�rv!�@%�<~�N�m�:��`*��0g	���ChjNl���Y��'}�h�wh����;��H�=�|�o{"�N��bA�	�xGroL��R�0���_���Y*���X�(�D`�F"M�g�A�\,�
M�q��h	�*�e���玴����,�y��]�2iGE�4�3o���`��
�3����xC ^S���[DO�2��O+F#S��q�A�^F��G҃�aE�7�f�!�����\@�Y�K�a�V�8�"�'�8��"��4�/ښ����,75� �)�^/��n��<-!1�-�Ę���* �]��U��q��Iv���E�Le8���T�@x�Z��}���K��,Wn���]7L�K�~sU
a��M��{��}Y����t��$m]��&긘s�������DJYJE0QΚƐ�4`oy;�)D=��0J��ͽ<�WY"�m��,�1}.��i��Z�1?�n��s9x������pI�
��"�`'����&EE��s��~�'ܩ1��b��0�7)���ͫ����ъpD7Z%pJ��C�*����a�$A_-5HXAe��;8+�:��W���ƒ���f���p�	F��-�tm�XF?
� ŦX�� *kH�v�����-�N�uX��D!̯n�H�d&ބo�IB�0��&���F�:?����w-��(�=]��Y?"��ъiVv�o*f�lfA�:�K�=Z�B-
����*�dGQ,�sW�v����bS��[yI{��/�3s�����$TAަ+�er����fufx��DPj<m&i=����D�܍�Z݀�z�2����A�j4 ���K�N9�M�@�����ˠ3���b��ϙjP�=h�%�H���i�O�����u�����N�cI�/�?�߬�]�v~�|������QӪK�aX ���ä��bO�:�0G���-ۡzF���u�3W�;4���09*G��s��?�i��a�!�6�������;\"a9n�^����@%!%y��S�C��Y�C�u�L�u�p5bg%H<G@h��Q�Q7�j�i���G|���u�2K�c�+nU�w���/����|�`H�9��L�wˁ��Y^�?�˾�;��II�Q��AfWt��M]���h���Gv���}:=j�L�M;A�Zi��x�Z�X�oT��-���K`������G<\>�,��x;A�!=�a}�@��+�������"��17�vZ��=�v�J��P��1���}��箚��+��^S^k���Z�a�L�xMeϴB0�D�k�$`��� ����ͫ?�`��R��'�d��?8g�#hA^��Yl�'y��r���R�hzĺ��Zc5wAIR��;.	wge��!7M�ea��܃����'{�up���Fۄ�B���k1�R�x�˂����#ٲµ�p�0<�%1?Ǎ�܁�q��2%=��TV�;�b*��+����)���4��ۚ���hqz�wǛH��Њ/ת�Ǭ��������
\?�T�=��x[CQ4%n
c��9���K*���S�c��C�#�
H�9���}�%��&
u~u��IC㿟U��l��h�{�OgF��`9DJ,o`��$�Ɛg9���$ �հ�̽9xI"̙�F�ۀ������z�3Ȼn"sÊ�#�ܝ@Bθb.A[�`'S%���U������c���%ʘ�ũs4�<׻���GSCw������F��x�����o]���e���Q�[���mM4��(͕�r�BS�h�u�����Q\@�*�`�	�F�Êێz�a6��T<�M�P�����U1��$�f�j$��A�"l)
s�1����n'�[������Ԍ������&�6�U��T��L�C�ə�M�̿�Eط%�|]�f��m�P�x��+51���M.>���T�R��7�:�۬� �>x��)Yd�<a�c�5M�c��X0k��zp#8*'zC��-�h.#d�,�7jj ?'GD�����t=b@�w6�Ѥ������'�]v7�	)��a�[J xU�B��S���a�?&�z~Oa��{�fzjAb�R>s����ye���r+�����>vI�������5�W04������u�@ED��܊��p9��I8��	}Kd�*,�"����HY����%�3MY���U�7vls�c:"��)�H�aO_
��gy P)̒�8ln#]i�=v���L����b1�Y� .�fA>����:vh�.\%��`w��Fg�F� #�� !��S���Ԙ����팔`���N���&���G��M�c���{�MCo�H�H{���ŕ7R�4>��w�k�&'!�>	��E;d�� _�S�[��O��$"BP���(�"�o	�&
Oi?>G�,��Q���V�£�t0��ԑe2L�IYx��r��hшnN�,~�ϡ� yl{#�w@�����ä�6w ���T��\�*ʮ�l���W��������B�\�r��L�U���^�];�@�/�c������!,/� 's�'<�.��:��(��)�Sτ�K7��Z_1I,� ����e�_���eN�l��?x��3C��*�B+��(����o���{��,���,�ou�3�+}�-D��eC��ӧ1������ϰ�݆��M�9[��HF��S6+����n͟\q�����`Ʊkj�|1<��a�T<g6�ex�l,��^
]@��_1E�>��dg�y����jB���x��k./�)6d�ly~+}mP0�8��IsQ`�f S*E��~���s}:R��r@g�cI�V+^���SA��:c�f^_����IP*\5�T�+���rE�K���'��� ����ɑkh�E�a��J�L����9S"�ϒ�L1�$U��O��k�~5ɂ�4�!~����k�0��H�*}�?G$g���kY�����HV�ܤ��tw���YiV���0Ҷ�iQ���n� I�8�u}��N�����ݼ7Ch���������|ԱU�<��,�֐"�I�Ҳ�f^:x��D%Dŏ'�d�ơY� P��kv=�9�j���`�t|%]�
&2�Eg帩V>[���9�[I F�Q?&�+�)�0��A��
O��3�K��9�叺��.�0��&����� �h$�9򲜱ꈋUrNwG���bR=T+(Q;��)(-�a�s~���-:Ϧ5��b�dN\R1��n�nx���8& �c�<G�e��|+|��)YɅ
a-Z�=;���p�J�{O�N��8��CT'�K���+��`bբ���J=�&%�r,�_��b��33q�f��A���+J�#'�\9�c#�x�����=P�YQ?��!^��܂V�]%��KG��+�<*-t�,3n��u�p����"����<��H��-��hk%��XkF��ڃ-d%8V�DlU*��},�)�W^b-W�	�p���(�����;V_Y� 	>2! ���S�0e��"����۹_C`a�/&}*� ��t�Hc��Q�Q9{` fm��:�JB��� �\�5�#SLœ�|�)B�[%�C���΅���>�!�R%���y4�Ѭu�}�-�yE��� p~F -cf<	���u��s���b��zu�[ȺA�,��{m�Ð��e0�(O�_�M�7���s��ۊ^��2�?�V�|�BaZ��iSD�����7�@�bgQޒ��S� Tkۍo���"_|���|5kG���=�qPr�T%���ȇx]O��F��0E���jL�܏���C��']��=C�{>Z���E�h-!���xC����'��x������
4����=f/����������a�����7���'f�'ʥK�'0,���q����v�I�SW4��� hV�X����O�!շCN�
�N����wt����}���hvK���h��k6��o\>�fA���~�q��ȩ� � &R��bs&�>�v��zE����6��W��7������QL��tB�}q0|��-�]dM.M�G�d;Щ�>|HE����Z3&B��{"S��DOʔ�?RIN�;a�uM\�9�Z��y��h�N�I��8`d�l�����k�k�Y���;�g�
LߪAj�@S{�ߤ���ö��rAO�iS���1��0�P�h]LB7�����h�_I�O�8��ۯ�ߡ�(f��Zc �d�E���8�D�s���X�ƵG7��&�m�
8�\x�ȁ����� ��o��~a���n����0�g#�1?�y�5=�c�My����xT��yŉ���l.>,o'�
M�9�Lݗ���Y�8��9%?9Y��,V�6Oy�������n�,쇷�_����/�L6��޶ȹ�T��~��7�n�ޗ֍+��<{�Ao=�o$�n��e%>� �ҵr{��M�]�w�%Et��/��UH��=S�Xt\���B�$���� �:0|�C�Du��H�g���rv����*�c=g8���0�5~�f]��K�t|�tl��)�CF�2�U��(�4{�"�X�3����E<wl./�D�#����ޙ��'�<�����.�X�m��D{�Ǹ���]ɜ�?��
~��7s���¡���&�Zc��^7�-HSYJo#�@��A�������],Q��^v�:��? 5�+u/�Y�}/:�?k��	�?��}]�|*�/@}>ձg��V�{�GC�,�-~�x���p�b�l�[��CܼFɀ5�x��v�7�@,rjAz����k�D�V�|�!��S�{`��HsX|�{Y��U�vM�p�w�d�����nH&/�$qX7��d" �3G2C��ۊ|�P#�Nu �$��.�3���i��s�V�3�����x}i�n�?wj�0�=�d?�	�t��F���G��?�TP�z��cEo�.�?.��~M�����Kw4|����(Ce�D�m�b��(��^Ň7Gn�V�Fv�ڳZ�}���ں�:Pr���κ��2Va���O�f�04`�Si|����h\x��<9R��Ԯ2��5��@Gk>ܮ&�T�R$��F��d-�U���`[�Ak*�����fY\��Uն�3����&C�T;���WI��vݠF�֨��QA��Q0B[ź�e�J�����z�t�C'2o�T�A蝕��'
vq���*�q	k��&L�h���J�:��_��9´�+��w���n&�q�߁Z��Yk�~{YfB�9 �~E.l."���l�*}����ܚ*-���AuD�.��GpQ��*K��X0�':G����FYf�}5��#.��Q&$�oS���~)�����%���7��z�Dڬz.Z�'�ԁ���b3�-�}h't�~R%�s�ח�����		Y]}G�#�⍖q�8�"i��^����toqer��,К�/Nߕ�s�H��&��]�ף�,F�cʛ �A�C� �"�ˤ��d�����f-�yTJ+fg<+�C���aP吮���d����9_���m	}�q�;k f���1����K�G��ȵr�~\o��R�{A=\�3�ȹT,�˷>�J�3�qnw���~?�����'���q)Y���;�F�Tѩ�?IC�F��+d�'�p=��5��Y| 8B�;����yC���$Bx2ͷ��P�8�ؖek�/�)E_��	�s$�q��i���&6l]
�鍹�HJ^����a�c�AN�ǩ#ڄ�%��kWԗM�,�9�"�If�]�<����o��"��m69pb���h�)�ϕ!BfJ0�JC��J���V�*ymq�ڶxuqv)���\�_�+us���eB�\���IB���
�tU����;k?"���\ג���f�P[���C�wD��L������S𼼝�� ��a�����n������v�D[F':�)E�=-ɥ��U$�p�aXx�#�?_5B�9)o�D�< ���~	:�fA>&_ˣ
މ�h��tH�	�e�@_�L`�缤�1Yz��4�NPEӗu4[�A!�G?p�Bv�Ӥ��?�"�pU��׌�#�^v�O���	s��C�S"�	���¬�>���)/wm�R+����rr�#y��{�Е2\���r*��%4��PפY:�9���\A%(�M�$�2��.{j����Dc.�Z�b<�fbo�*v%H�j�G_r��5+[p��� ��?Y`��|;�U-���Oa�O@�5��[��� d�����?f�|=zu�(��-�W�Ոb��I�0�OTL-�!����l���+	����fi�r@u�S��Oo kJp@�ӧ�MMْ�\��c��:�����+��4a<����R�%3p� R�1�4�� X�?�''�������'�����6�w��	,!�m�q���'�ID���kÓw��DXCH��u>~y�)���R6ES�$}?�+�5�"�T2Gu!�̸G�h��K?��78'��j���Z����>�ݯ�^�2g�C��-�X�	<z���s�eN�(&��\Щp��p�\`����+��a"HU �kz'O�4s��(3�m7����⼱��_6�ˑ���N�ڪN�8�4�Pծ�Y*J���7���}򱹕�a\HjgE>�o�b�����^�� (j���rb�o�9��tJ��B�iΓ��O9�,o��_s=��{��}k�s���4,��1Nݯ �Ce
F]c���U2^�Ԑ����]��(?At��r��t܊�xT��h �� �7�h4�]@�>���`Yk�s%��F��l�� mq��.-���2��؂�;f�By@\;�h����j3t���pE���n�~��ڲ8ղ�����.7�Mhuؒ�w@�ӱ�$Ր�W�����KS�e=�@[L�+��F04�e��L���n�,�8ڝ�u{W�d�x���˼c�?���	�L̻QB�wrt�Z��	�%�"YS��C��6���%6%{E�1~���(�8�"��9u����U�f֏�:����r�ὐ���� ��}nGWߗJ7�)�zA�	���8&�����Ԋ��H`�*����A��NL����-�솉~��n�+�؅��;�;�W���S�B��q������	�%��3�)T����1*0y��L_H��<<��gk�2x�S���|o�91��+�:�qf+q�H��}��v��5ʼ���DVbj�R�j�f��S��v�q�#_k,Z��J�� ��bA6�_�P6��p���n6�q�7p~]F�{�I瓷u��#�~�,WP.�:k^N%/��Q�Ƅ�3�d
�9��o��,l��mM����o.�B�z�H�>��#�?�-��t���Kd4����GK&)�ð�^�û��qe�D�G&���[�ޣ������)���$l�F"�5��D�s���d�6��
��1I��{� C����{K�u�ɭ��E ]����tX}o=Z���U�-:T�C��U�&�ţ>\�h5��@�eΕ�t�a	���>4/$k��+�Z�\\T|0���C>�]�g��B�{mf��&qx�{���s����
�dW#ɰ7�xp}Sl?���[��|.j��[ׂ�h�>u
ȏ�.��I�T!��e���H�NCu��&���M�U�h&�t���
 1 'L�>���y,����h�菃�m����o�5�X_�0����E��)�B���,@p=��7�7����`�l�4'�n{_��H�Q��B�<�e[%s �x�Dq
�&�t�ԗ�,�X3iS|��.#�8#��Q�Ӽb��$e�⇸�D�"by1��B�̐Y;���u�M#��(�9
�&�9�M"S064�o�]J05�xD{�Tӳ@�u/	�IHt��BwjgI�n�F�B2�����;�f�P_���VQTmM�}_&oi���Z���4���?��`��KF}�8�u���\�`��|�N�>�",j��Cʫ��T�k��>C5����8u�*��e���M��`	�9��O;�#��U�H/�����uxDu1�*n��$���l!#�;n���C�I�����7�Ӷ����	+����`�K��6�?�TJ��I#���Ӏ��\�e���ϋM�P�5�[-�5����N�����U�]�L`onA�cKQ�LF�O�n��raazѶ �a��L� ը��ά����"d��)�Ȟ�6֑Rǎ�ֶI<�@�Y�慠�%
!0�f�ȫL*{��e� Z|sL+��iһ[ mf\�D)��pH�O�kbJ�|0{��i�Q ?��Gx+�iB����Ѕ4ǻ���Ǽ"�2)��y�󛹡��_j�hT�%Cl[�R	4������+�`��7~�[�9�X����~��5Lqk��lY�2�|���;��Ƈ���v�!����7!h�(\&/Ġ�Vo>#�Bҫ����W%�;���r˓:D�{������$c��C���z�`����2(%��
o#����8y׻r����T@��t$TNK�J̓b�M�~>��d��׼eo6���)�t4�C�N�8[>��(��jǂX��i0Hq�L�Z:��i=�0��2��`
|���P��w/T���S��I���I���
V��z�EG���R��o���̇,��O�L{ 3��f3޽_��|��D#ʷ��}&�*�w��&� ��F���H��Pz�3Y�3_oj�u	�o�+;XL�H`o�mL|�&�`�d\%���rj�-�����Xç4aZ�֒�R�"�L��c�]�Q$`B���R��Ù���q��G"h*n�o0M��&=c��ڱ5کKt��oq��q���zC��Қ��t�if����`�'�
��i�(�[މ�ͱ�G���0�$���]ӽP��'F߫e�7���W��G6��� ϬlwZ�l�ض���?�~
v}���F	z]΂"OS����������R����'�TPg-�KүX�C�%��Gۮ����+#zh���&Bܹ��g}�I5�
���곍��[(�ky��qh�sr�RjAHC�۵�k�Be ��O��D��0�0��t��tBp���f6T.I
[l����mD�cV�
8d����ya
�!u���[��Ɋ}�7a���9�p������o]\��}ᑵI��}-����dJ!�<�,!�&q���TkvOHE�c�,�7��y�����4 ���NHԢ֟]���P�!��X� H�N	#���"�YÍh�ƵZ�����i�%��en3��@�b'������V$�XE�6ƸvKJj685Xh�p�����:p%�d0ltC��k����:)ɥ/yPI��%x:�re*��@�O�P�;$����8�
����A�S��Σʫ˻-Q��9~4������n�X���3����\WGx=�.�h2�)���i+�΁�L�=0�z���-X���8��曍���p����e��,"�u�[(���)ک�Ca\r�������D�s2��O�ڜ�,>���̚_�a懬v�1 ����R��MG�;���Lh:VuGz�x�P�!����Ֆj·lZ��>�2���l�s> M?������,�zn�;� TGn����2���`f�nI�)������Fq�����s?㼊���f�1��{���5�����mp����h�D"�Ny轺R��R?��Ju	��C�%�I�����dZȂ0�$��%��@D`y;��S�ϚM��y��_Kb`?y���q��J�]������X����OF����Ҭ���[��� @Ტ$�%|Ug@�p������-�ؚ��U��B�� 7�x k��P��\�Ȃ� �4��HzN�:7%��j����`iyKjE���5��T����&���0��޲!��8Iԭ��� ^r���M:cf�U'���᝾��DeP�QD��%_'�w���F\,C�?<yF��@�>���Iq���]���]��=j�} B�g���t����R�i���I����cҡ���E������ה�i@�E��)z3*��
\�W#�NƙZr����z���O��f_S�N���I?m�ZN�ׅ�&D�G�09��|w������PN&��I��9k��\m�"V����0i�`�B趹����4��o��!��`쭓:��J�tk�oT��
V�1���'D�����$ȷ��e~I��^1E�k/Q����s0ϐ�ɏ�!'*�?���e��s�Ls45X"��@��������𫍻B%7�f��ݴÏ�q �J��C��ĐhU�������<��mM���=]�"b�v[�e#;�iR��Hrel+�_�- 	f���Z��� �p�K���Pb�R�4���#���n��t������T�*>��}ۑs�e��e����W^a�ܴ�^�?�����s�`�F)��Fp��e� OA����گ��m�?k����Ht�7�f�z�}��9�SG��x�&���ms���a��
����<�2M�����ϓc�-��3]�GʝNٍkp�ݜ���OI#����H�z�eZK��ܐ6'���L���۞�X>�7 �`9X��+�}C��
\����]�0ty�~:Y<����yI}����P�w��|-k�(�Dąq�����>��[�n�}�f343�[ƀ����S�)�m�/�!�Px�+�7E�G�$�,�yM pe
���gic�Z]���?�Vw�-ك��ƫ ���7r�?��tL<���S	H�'�9k�҄әB2X�57����}HwU�N�O�� �ȳ�Ii��DE�5�#����U��w7N����k��P#�z*� �#�%��h�+.'��7=�ʦWY!`-/ӿ��/�K����N�3{U���t���� aP\A�~�LN�),8���ed�l�|�	Ir��)}�~�FІ�q׈�sK�Q�a�B���d��nq��o�cwZO�:q�(�S�/���+��7��>�9τ�1��0>����E2,(l�M�迍��|,((�;�3đ�zY4�*Y7X?e�R����9���?Q���{�<'�s����pS>�a�~o	pq�9���-{(��bN�HHD���)�V\S�h �Ō�y��j�Ƞ�P�!��ݨ;�� �#�RtMͨ�w�D�H�s���3:���kQ�ᄳRu�?�!*��n���඾ҭ[o �Va?Z����T�͚���ۘ����T�\ܑ^t[���p��DS�.o~����X�ZA[QH�E�8\��D�)��e��T�jR���߅�v�ԋ����>��E�v��+<��ۏ��_�`JF����r&3�$�0�::> R�9���:���G\A[�f��y�|}0���k�MJ���uu-y�:�T�L���	zv6 /���UVg�ju�R�fgAtLѓ�h��w����n�_-���Z)"�v옖��ER$BX}A��L;\���LY�[M��9��s̅c�$mc��P8��������Y��~MI��/���
-�_` �(Ui�l\8�]+4�*>8!r��`	����S�
rH�E�x��-�bf5�i���Mt^ʭ�Vy� \l��o$j�[L��5f���gO��-���~˃y�����8|�_)�����L����.�%����,�/9q��n��wp[��t)o���!;�	7��O�r2Yh͸wTP3�`�n���䬂�8�3B;\�,)X�l��ݙS*�����t`�倯�
�R���DE9��h�MH�,m�����T�V����B�E�m�7��o�<���T�m�6V�!�S�/�G�*��哰�B��/(���2]W.�o ��k��P�q:�y�03/�/a��p�D5�?5Gd4 L���tE����M��F��n����U�rp�v��A0�(̾!��U�NB���Ό�x�-��C�p-��=���C��Y/����s��(�ቺ���d�8w��{��,�������K���{�=_k9,6>�����XK����W#pR�X����D�,BK���>ܿ<c���.����MmއKnb�D>`Ƽ
M1��=sg��мc�^K�/���8���1=� u�5[Χr���y���z���fQ�'2MqS���1]N<R2p/����e���7Ng��)���-ӦF��5	N��.�儒�҇�4>��fY��nG󟦸�zh��<��C����AO�3[P�_��y�)��X�`F-����D;�{%�1� W���g�a�AW��x"dg%铱6��,I�Ѝz\��6�1oD�_%�B�Ƃ�����.o(T:'��9{E�;r�P��B�� ���O��B��q��NVE�]���Q�(1�j,g�Lc�kC��=U;�te(o�*s��-G�,?�?uV����s��x���DN~��F�qP��7�dh�.:t+�C�����s���oL����GD/�SX` �nP	 A)Yk�C���C��CE�������E��N'��6"L�皊�-��0?�Q�J�Hi.3ǌ�sB�5D%�U	{-�n�&��}���@���+I�2&�F(X�����P�0.=���M��L��]��[4�n���Lͧ*�P���a�`���*7�xe较)������b{�.f�%'i@G;��D�"9\��z��}/i�L�z"��)�)1�!��B�r�����K�R��Y6��m��,��"ˉ���aZf1��)e�V�d6�8O��R�[�.�@[y#�f����Ƥ�g�4ٕ�0"$�]���Ͼ6��2��V�/3����;�N���3V��Ջ��^rd�O�$�:��5j�I���,���n؅`�׆=�+4��W#8~�VpB�BZ�dPj�Q�>6�,���`X�	~d��1�6E3��b�m�(y�g��^�^�8�=�C�:��o��	��uڳ�D���-B�rF���Ϛ�$���1��jG�m^�R���T)��o3 ����_��Ry��%KX��1��Kc8|���yJi�%-8���u����Ty�ert�Z!�vH|>������O�xXG?nR8j[E��D roFW�G����B�k�_�1ʅ�"X�*d���Y�wGА%�l��Bt�F�s�6�T��0r.��C�D��|5'j𛊫�����a&��B�P��`�փ"N s(�F#@ ��T�j��l>�8�6e{���h!���_��;b���ʂ=ýYG"��z>w��_�2Mr��Z��Ⱥ���m�Z�˸鬠�+ӝv���ߩ��ZP5sn�^i=������BG7.=TR�g��\�l���S.��d�x�J[YZ6�%Q[�D*�%���j��:�"�.����#�k��ݹ����������$"35����H
�PP֮�Z���a��� f<@��C/��TvA.V~�+b���(�R;rB�̥0�T<&~?EĮ͎�����JI��Gϫpg� ~���3<S��<�z�mW7�,oi/Ur���	��L&:P�����<�� �9ĵ�Dr4�麽]ɲިl�h[�>%])D�n�8�����O�&�|ϧ���@0�}���ޱK���8�*���-]�_C����,=�$��[��ƈ�X
�8ZDæ�3(���ޔ����5�C�Jw5�r��>�[jɜO���޵���Pl[�_����
����L�Fy����2�M���P�۸@?��ځ���B���_�S=-�ӦQ��.��p.u���u��9H�_Q���aQ(a[#�DG�<��1��p���r'�h+������$y5��#:	 �nv�K��es���Qjt�+�p%�-:��[]ڂ��Bwg�iC�����������,�D�4L]���X�K;MZ������m���I3Q�����A:�eMX�ye���8%�1�g���i}_z��G��i���ꥑ�Ͼ����P.D�29��z��⒊��Ԫ}����;Ds�=�4%QͳUGOZFb1�YU T^��#���^�oy�:�����4z,�nꮬA+� �W�z-�bVg��@�͖��=ʥR�Y�,� ���;��W.��3���u/��D=M|�Y�a+T�o\��(S�v;Fo=�[���ԩwE� ���0�������`�f�8YI5���n�M���e��6:�\��{���J
��Zq�I��d����WVuZ�T�6TK�,��3'o��F�_�04
KD�R�[T�H����4��E=֦QUAz�D�U�pPˏ+{_ݮw��ky}�٣��� .�)��HKᲞ���+gJT���U�U��@�>�t�[[%n��#�R����Ap��8��_��T�{�Wj�	��:ժ��B���!O �j�l���{�s��#jq�VɈ�m�I���_��M,wP��(��%L���@�[��S��cz4�5s5S�?��[q�|���L�|��ƬF!��Q�� ΡL��XyyL��1��ъ��ă�z�bT�h�gv����Y�p���� �yJ[]O�<&k&�#U����F3�H��fkګ$����0��oW�Ş}�^lP�ӯ��k}Zuнt@ �k�6�́HQg! �Ł����k����o7X�[��Ŵ:�}ྉ�,���3e����ݦ��d��,�Z�5oC�.$Iˁ��A��r��C.�����T��a�<��Ss��l����U�<��5��#Q��;4ĒH%+��2,�\�h3��)���]�C���R�X���h`ʇ�Z�h8�2C��;x������ʡ	��*$<E�gF�i���W�^b<��ms?���D�L���=eV��^_ ����"?�+ a�mR�I�1L�Z�����_�m�b����T Q��Ÿ�Ҫ%z~n�!p�Vd_j)���]�/���7��q"T�C�7�5�[��P�&2�ǟH�n�䅥W����o�dGzo͛u��=����(��wCZV)���+v���ة������3/N��L<�̷~9��+�_�0&���Q֖��o9C�Mj>§Gh�w�cNT�q�zj:}��kn=�J��O����|$���]��D�!F�1u�]��wlW�����3�e�A���u��W;�5�����\�-��0��qt[�(���J�·��Z�b�����'�J�H��S��9����.B�*�$�_�3`҈\I�OP�{�w����N4������I�ִa�h�:������&�q{����E����_]͛�x�D��xܰ� ���(�ĩ����R�1M������i@��`�L[K������~8"E���!�]�8m.��A�ꉰ�殖X7`H�q�=zw  ��Bt:�(�	��虜Eϯ�A�R�[���.�C5}�A�� ol�����s�S��X�w7��=�ˆ7�/��b>�x%Uj��쁛�m�h�4j��?D�.'�HoI�y1R�]jyb"t�3���6�HԤx���yZ���n�*��ڿ��%�ý��=]$�N��uo��<$�ǦY9�au��v������C6��),�Ƥ]~]����
Q}�����k��=��e�	��@�E�qC9���Z��\8[1�*S�C%աsC,T,׳���J��1B�۱�C�'\�bi�GǱ���^O-�I'Ԫ#�{�AC���	?�r�s�v�(���Æ(PB`San���]����~h,kÌ�����w��w3�S�H���w<�ٹU�JD9���f �Yf���A��~��4�>7��uF�޵Ų�V��;|z��2��4���'q�T���V�u9A����W�El)�kZ΁MrNRG�^OZg*�c�.g<� lj��6:�H�8�m{FN���_�����r��\p\Ç"-xԘhє �1mL�E�x���6��_ǝ����>�ze��}9�d��nRzj������"H?���	U2��Y`�1�5y.:�Ε�!fw&;�.s���/?X\��I����f��G�v��1��r����<6�T9H�Z�o4U�Ǎz������&u��
Z���[��^r/ �m�(CߣZ�[�>�#�'��3�8����`r.���'"�Z�������[;_��?Q��a葷�~�8�.�B��!��>e!��Gh��fЂ�����b-5B��am<l7���A%F2��P�U���-���qs�H��o��ݨ�Y�e-r>Ŗ�^[���y�-L���O&���X�ĩD��;��I��5hxB6^��&[3g\������^��������}��9u�m�A{r�s)���HԖ�o@k]�(�[H_O$�Q���^)4�M]n-+���&H׿;�O,;�n>Jޙ�
��Djn]��?G��]��j�R�Me5��m�_�Ti��yn ��V�sK!��j�=�9�L�+i�a���Bc?��9�6Ђge(�A3D��e��34���y!A���v�P��hT2|aX�*[$ ���5�o����=-�����޻��W�$� _I ����G�2�4~;����8M���yao(��8~k��8Qq��/h�'|�t}@���[^}3�޳a�#�_T����'���;�?�3�������q�����[$���vQB�0���jڢ� ��ݿ-|�we`���&t��c%8VN\�ڎ��ӕI'&��Ue��`�d��ıV�f�Bs~M?\ ��w>�(p�&%ps̕��oTh�&��,��	��KP�BPk_��ˬ���eb�����v����#*!���S�}K���HV��g�1�lq�W�(����8�Sl�IdBbW���a"ӝL�d���M<M�@�t��pL/.V�Pͳf�-��4��~��#��2���Z��#��e��T��WX@������{Dv�	A��)(�j��*|JIq�hBľ���;�)�̄���}.����� {��COt��}��������'��/Q��c��|�x��%�9���(����ٴ�ʦ�������Ƴ�%V���c����`��=T�����!WG]�9w_H��*dc�Gub�_K��:ݜ�0��`j��"ߡ ����R+X��h�zkt�n\Oသ<���1?�Lc����$��:���=�
�G�� [XA��4wځ�(���~~���&�b�{��%����W���_�j%B4c n��r�[׽/	����	s#kO'�n���+�����p29�M��R�\�dPtN��Ъf�EZP������\s�X� SZ��aP4������%�ufoI�?�������|HyC������^,d����;I���"���h|����6��0�����A�C����j!�es���ߤ-1�(�$n�kû��Y���,#)���pu�H����j��!d�F�)HrIT&u�{���mk������t�\��_Oi�K��W}����@;K��)�k�N�I�wSH)�B1T��V����oXѪ�,������c��\9;��oȒ�F>�Vj�?&�iM˜��{�Z���M�� �7���9}Btٵ��}��լQ�8�/ʢ�[�:�H�t�!I���BF�32>A�S�W�&�Eӥ�V�wP����_��RxA���;�g�q��fn�ۛ��0�1�����@.L�����e�i�	� ��*�F���,`���*c���m���A�AB��Ǥ&��6�R>bPZ.�g��Nm�ߣ�*,�e ��2�HqAd�'K|�DQ+���Tf�,�Q�� �b�6#,^?��Ϛ'��`��=���d'�M۾r� ����F"⿡Ք>���ݾ_��غ�����W.��mB������~�D�9t��E�PŅ���?�� <������"`��#��((](�A���pxy�Hݨ�1���x�7-�WQW�[�A�"y�f{���`t3�:�����6I�F���*�h�	�Q3K�������^$ La�0P�J��1�B��%�ݷ18� oә��2��=_&^�r�AJ�	H��g��xu3*߸��.��HwI��F{�1��ծF��Cˀ�*�5\���N�������)��A��n�H�ڭ�$?N!�GCx�"���;8���j5�ŹMz"R�<�zޚ��A��0-uo����+vB�!Ynz_��ߢ�ض
]mv0�-A��s���<,��Ŝ�����^�vZ%�S���:"��ۺ���B웘�\�ND�Q.[G!	܉aCe�E�u%f\��.��h�U���8���,��E+
�/��;����B1�{�Y!�
�]]�� �d��3���"P5hy��Y��N�������83uC��٣!��r�z|}�XZ�_�V����ܮ��܋K��ߦ�Ħ��>_d�>L5�����Y� �KMk�! �<Pvx�g����<G�8�,-�tr-Gz�7�����<Q����{��qc�iZ�`6�/t���8���D�D*Fclf�4�"X��LslE�ҹ�}(�Y)�����c�� D�y�X?At�����a�ǥ����6\�Pq�e�zO�N��^h, ���(6���5�vXU�"����� h�Һ"�El�;f���]��%s���s.m��t�A�Qg�t��^#_>)ۋ��iD�M�ɺ�J�M�m��̇.p�s�nx��X��Ԡ{��-%-���N����gA��}u=z"|\�lF`�L	�W���;
��������sp:.S�Vr�3��?��bs׼�ɢ�4�D��8��Pjy�����@�_Z����k��vܪ�Y&����� ��2�y9�ާ���_�[��ϫ%��Jnu�E� ���|,�U�������P2S�-؟�W1���VݮH՘q���?�;��w�7��\�<mS(������2�f���
5�6��I�A<9��iFy=&u6"�&�Z&�;���Hr%y7~���XЋDe������hQ�H��yA�ZW��vw�3�'b)�@� �ս�Zo�t���hG=%��z�jY���⎊��q�3�Fڥ�f�-�����A�_e<��e��T������X�|r߸oL�dT��¶w�7a��Cp�!!MOH�ё����q�	 ��p8��F0sE��N�H���W`[sȞ�NӅ#luLȟz�`���Sb�;Ҡ��W�����WE]�0�j���#l�e��=�^���T�}9��Pe�Ǘd"T_�{f��S��M¹zNT��Z�O`�������G,��	�UOU4��Axp��B,Ȍ�s�8@Y���ְ��DmD��_������h�,I�nsya=���S�ϳZ�\[S]����;�e���t��Ɓ�UC��G �;w �:]�@>��A�@.�^D�1���c=�٢�L8�_��taB%��\:'��OT6�� �|�yz�`��$�iS�{\�H���d�����3�{}X�	-܅L� �b�$1&_�$��d�"8��xTݔgKC�����폢7��� 2X9�s������������p���:�o��/VS�q
I�' ��a��)rJs@����L�p����p�\�AK�K8f�#��]uwnye7�� ���GЂ&��E
P�v%%�A��b�j���L��ZKFP>ܓ��q]�����&^l�K�[Oa?0E�H[�09��6`��C��q�ay�Ɂ�7�~���8���!f����o�h�3%uP�;�YhJ���xD��oW��=-�[A,��YGY[.���~�<|�#���#�<(J���͌ Z��F������y��5*�Ӓ����^��h�7��Ғ��L�Q��5��%�Hb���p�t�#[�*�[�4����PD4qt_$���DHh
��
��C������>��=0r.ۨ����+���=L޷��;�Ô���(��~��_���U���z�K���ΐ`c\��9	�c}t�>�!?V+ �vX�{�J��M@��Ԣ��0O�NRN�@n����`�W
L�=XqrǃϢ'�p��1k���v^ /�t�b#��I��4B���4�1�V�����Xق�?Ƹ�/}��f]�(:���m��e�*��鍱�&�q�0o��χnn<w�n��9k�s��@4��S3/TNy:�g�<��9
Iސ���ӧ�����\X��8㲎Gf���M.;����1
���j`���(���4~J��W8��(N��{ �o6�8S�O	-Y�Ӈ@���26I���ܝ��0��5�p߉3��ޔ5 �p�$�
Ě�~ � p��- |��Z^�!7��h����׿L�sQҷ�(��b���JO=F�R��ˬ�Bz
?a�o|� w^aK��_f�x1-���4�	{�����Y���1�a��i�+�z0܊%Pn�S��P��p�9�+bkb Ҧʃ��� �8���Tu��L� �nN�O�hAA��ӻ���5ɚ�t+�6�[���@�K=�J��ʩ�q��Բ�BK��j��`��/[�
��_�~���g
(��H�#:3iTK��Ѵ0��)I��?���&h(l��#m�$"b���3_߮|�W[�+- 	��֭OԢXN�ޒ��cA��ھx�C6l�?7�*�.�dh�g%�j˃�=J�E��MɌ(��^i�9Ϭb�X�A� NC�7~��Oܤ�R�^nH�̢#?��B<F�L��o�����m<��pl�p���V��Z��$o4H�����U���]���V��zC � Co���4T�f��(G��:SjDTeI@NS�#��mH�;�w�{�Gu�]��CB�ԋ�'��3T�?|_�7	��B5�L����=u�|��=�h���� �����>��w��6���q��	�� �dJ��T+B�6�(����ʿl�	P*����8b�;�!�u�p/f^���/�R
�r���;�*>���z|��8��EWύ�o_��V����A�ti�3�rg��;�3������iT��Hб��9h�0ef%��tiU��\7���؅T^^���)����)���ގh��T������S7��Ｋ�/��ɫep���LvX���&s�����g�eӛѨ�%����n�l���������{I,^�R���f#|�3�;c)E6%�
�WKg��?�՜*Pj )(���Y���=��E��K�wߟ�h 5�B��=��}V*�`�)�k�K]�Ēz�x(���-��{PV7'hG��6�ӊr���H'$�F���wg��q�O��,��k���I���bZ9B���d�Jf���g�X���ι[������X� ��Y�q�af�;�R�u��97�%<a;9�����>!��z�4 w��"Y(����jN��G7H4��F[��D��<I�B�p; ���U�µ���b��D�3�K��FG0�'�$�aMA2����	�`0�- ����>ep"�x�F1�t�
� �T\nЭ�e��p����BJvƍ{�.���j���m�����K�>�Jp�rYƍ<z��s�J��XC�SlR�15��p���*�v�a�7?�t�Y�]�������f	���R:BE�������y{��$�ȝBIl�¿�o���L��lb���h�5�f����z�Ʒ�QS�~����.�w��$�y��?�tlU�D�	�)���
\Lҥ�Xj�1J�:Pc>Wd(�m���86����±�^ы�	c�<�sE��B��)ÿ!�ؗ� K���<˱��{R�yk�Scm̨<%#��rZ62�/j���zY�9�^P,&�C����e�7��@����xn~|�J$��3��[�{C�;��� 曈w�=����B��%s�=mL�si�4=�0cD�B��v���^�����PN�
���D1�}����D���׻��Gǂ��Ӟ:Gom���_��O�1�q�:kO��JW��*u-4��Do~�3q0�a��Y}�����O�Y� 8���g��b�f��4 ���I�R���~
�',$�D@ޏ���'�</�Ǟ�]��d}BF��R���v������V���� E	烮`*�$�1��A���1�����g�c~6�鴷	6=?AKWC��b*ɯ�E���k���@���N���&V�V���;� ��
 u���X����f���pgw��y�:��7C�G�*?Fr�2D�Nxy ����L��f1"k˨L~px�H1ޛg�v=��-J�
w̺���HXNM b)��]���kB,�r��H(o�vN$}�x�+"SD�\�h l�t���Mć�"[j^U�]$P,aA�ڦT���mF�ن�(��BQ�B�KT�]�}�BΑ6��]g��~��u���%C����Oݸ=���*��؜�r�\���/5W�O�j8�-��ڸ��Y�ji�Of�"���Ε�y��U\������w�il#�}��*eM��T�zV��Ҟ���6c�Q�U��N^��n����lp�k�ڃ�a�4J����Y^d)���RD��o�|u��Y`��r�꓅%a��:={)���
P!����.��,��l�#��,��k�d�\��)�`���O�WX��#�=`ȫ����0TV
�o�D+��>��Z]@�3<L��=��`U ��(}�L�3[��B��S��x� �¢ �;}��+�>�б_f�Fث+w�N�t5w!��^�;��L�,��ⴈ8qM����^-e
07U��`H�7�mˁ����ǳ��4P7�],l�nl؉�7�!���$��ikr�ym�k������/��{,$<`�>��2�;��y���+���|��m��ͳ�e����5:�3N���5fp��D�Ta���n�� �S-��¡��2�Bc��d����=������
�2��y�.T�!;C�Ő��U'� P���lId�P���.�4�G�!���BԮ`�$΄��?"���UA�/��Շ@�˞�0��'В��ڶa&?�'i�.�������X�R����*����I�:�\�|�V�yv�{\Ǆ�1v�y�ꪅR�B� xSn�+�L(��(�<��G�^�. xO��>�2\\*�Jyr�g�#P�u���K\���S�}F���+Ԅ���x � �u;͸��X3�U"��sc2�w%Ξs�Cj"ꄩ���i��X��iU��A⫔t�Eo�2��5)��O�"]�j<���nK׼�q!��Uǫ`�M��=n����汪��%�6��>a�̬�F��)��ƹ�(.e<J� pI���߂W�d��(r����%���Wd�������X���f}����:r� Y;෴�)��޷�#�j	{��xV!����ۥ��S!\�U��������9���B��ۙ�<��T�Zs��"?h�@�W'2!(�I=��g��R]�dT�������ؘ�R��,�8����C3�O���ֳ^�y����{
��\w��F�����X�5���o���!1�ؤ�7m��`�N1̄���.| d*$đ����*��`H?}͡�T�*Kz��Q�L�J�����v�B���8��'q�9�����>�+�����NnT�nU����uۡZ�ag�-C��.j6q`}�E�,?�+*j{�� �0W2g��BSW�i�e��8ǐ4��m.�{�!��[;�&f;��⽅�gy���#x��a̢�.B/j�N��WX���Q��O�᳡��ѥqԕ5L��VQ7��������-,�Q�W���(c����6���tLj��jMś��̗ g]F^�'��n��c^V%v��|�.�+3M[��� 	Н>�`W�
�o�F��ݭ/&9�[�'ni��#/�P��HW��6���<���S�s�6QGc�ٮ���X����LyCBY�{Lx�v�� H'uf�]g\���(�|�2�j�d���E�t�֋k8C����q9�scB�k�z#��ű��.d@��� �Cqx}�nܠ��0��9��˶h���� d��&yG�g����+�hR-�����"ߔC����a�I��{&���㕻ͤ��mX�U��WH^tZ|o(SC�[��Ǘn0��-��9��tNz ���}z��d���^F�j�:�u{��Wv��>����i^�Yg>&ٷ�'���6vy�|v`�6��$/�kn�2���ͣ��2@o[�������g+f>$-���t!U��TNdp>��tH����nİ��Q�@��	1����<m����Er ,Z��j�ӕ�j%v�M� �u(������+r8�Q�&�qb	E�9�����}�op�'��x*9؁�	q��wD�S��eg;˙ʹ�;?i�C-]f�&|��T4Eh�^�n�"a$#�t�-�����҆�WWr%;E{s�<�T����~C���}F|pv�7GVՅg�˫;배U�ԉ� <�&�����"��@'+ޝ��A��Ft��ߝ�%�?�d}���2Fi˒�$2'�}Lؙ�5)(kQo����:��{mX��ԁ����V!<��=R�����r�g�`F� �J��Mw5HwBU[������d���I�BX�p2f)��Z���u�ag�qSB4E��4�����S*�,Z-���׊4�쇏�V�}�RF$p�P����j�LI)XΕ������{�f�:�n�l����w�w蒍�Kv�
�������A�Rk�"�pJ�췈##G.<�R��
�5��1�����	�;���ƴ,v^^�wR��JwM]�û����4��j��M��fk�p=��x�}�q�����2ѕ�"D������ؓ9u;��)O�[p��� |͚!�֍F�bg�R���~^m8�D�y2"��ٍ�4K���d�&��/�@F��D�.a�G�����B�f�=��,�VzFӳs��I�psb�EJ_;L�d�l#`:W�7��8 ����머_y��ԃ������@@wP�E�%C���E�x�e��g����h�h]H�M
�a���$+�?�$;��8)ȹ�0<$�o>�\*���.A�A��H�U��UL@<����+���b�@�5�)��s�ʲIv�Q&/Z��!����.s��ʃ�]�jpV��zE��d�����[_�s�*0����4g<�����	[���
aS+#��m[ԖɅ���Y��'�N,���_�&)�ό�+Bw�[&�����I���xj5����(P���uz�D��c�e�c�B����@��_�`�	�Ƒ��o��[wp�d�����!W��HJ"��#sm�����`J�`�`y���C�3�w��'�Z��ܟ�������Y�`�wD�9J	�HA~ۙY��]����~�@��\p�Ӕ[��?I�&�Jv�,��R`7h�9���A�.k+�y��ypϩ^(�1$a��/��<1κƌ���2����Ku=�By�_�"�v�3�*����Bɍ�dw��0�(��K
֥7'�JsqD~эeڸ6:L��VpU~�.Y�ĈfF_ex���QV7ީ %���V<����:�{���c!�%�9��������؆�ʏ������(��o�|��ۆ<yq���z�M�䛨V�ْ{&������̐�pAu�Y{E�#pqi�w"v+��DAz�����S��`n���a�>0�ˋ/82�Ť��ܽZ?�\��T�XʳٵV�[��`Zޗ���g��p�â ��f$���4���j�e����~�|�Q�9-y�Ġ� ���Rg�L1���Hd�F�s>���b *�x��Z�~b´Oi�͓�#H\�}2�e� �ČāK!8�W�ȗ(�k�[_,M���֮!��b�G`��#̬�%,֒9�P(&�������:F4��&��G�U��>��JK�=�2�����6qﯼ�����c���hDZPY�;�t@��uvUċԨ��`�)�
�S�����9�_���Cg�H�z�m^�h0mN�<_zmW�a\���s��8�򍹤�=��;��\	ȣ��C�)�u��(�持m1	�~.Ez�k�����O�@G�����Ŧ}�Ǵ̱+���%EIZʔ�z������) OI��N���m�1�P� ��S� ��C=8��ok�w�Ht�jo�]*����pb���K$:u
~�Z+ �^E6�����Dt"@b��]��\�~tz+�"�O�zL���s��Ih�]�	,4WϊN��QT��g�dJ��vH�qޕ�={2A��1������(�К1�DB�(�V��*�%�Q?!�k�{ؕR8�x0����z���8��G�����B���f�+�Ǚ����u��ۜ>j��[[��w�県,ӷ�EO(C+�;)���@7Ŋ�*��8	ʂ��x�qUz�c�
�bh�5t!���O�W�<����ּ��y���zB��aT�������	!x�wŁ+!R���X��
&�RixV}K$S�!�գm�a�fdAQA6�����/�1��T
��/w�� vN6K7�~M��쏓� Iw��SZ]��MY̰=ޒ���Lr��p��;.x%���������?n�l�W��$,��8��B)^^��Q�6�co˖����##*��N�!� �R�*�����8
!/X��t���q��?�jb�d��?�e�������v� �.6�-H��b-7/�3���!*cjK!��Ҭ ;|�~��ei���ɬ8�8���!���s������WM�~����e:��b������}/u���Q�-~�Ӻ�^�{r�~�p[�D:*U�P&�R����Q� �i�K��1 �������C'��l��<��vhѴS��R4]��W�\qJ����[����z*ݷ�'F���-�M֗�jJ�7�dG�H��$~JX�zи�g���DÞ��̊���קN���V6��".�O:���PN�{jY��6I2��V���Q�9?@�.�5�?g�M�(�m��j������Z��i�a��i!H������]��%���/Hjs:�����	?��R�h�J� �6���	 bz�A���Y
0"ZO�*z�ra;�Ѡ+�a�D���:D�yw��?Қl_�R�_���@���֥2(�\��e� ��x%��v"?ϼ��8��?H��>�@�1Z!��F�S�԰3�W7Pj�3)ӎk6 �#��^&p�#[����@��沣@u ���k���$$��逡(��g�X�4Q�[p�c�߾҃-u!ׇ���N��46���`��?��.k�\c���vj>��G�Om����y�+������mϵ�E��)
@�=�i��%����W�Jď ����S*���H�6�"�ba������G<Z{w�wй<Q~�܃����\\Bmw۸�R��_����(�$̜?֓��C���"��?k����/� <~�{;������'���,�?���G���E�d8r����FԈfoz�Q��	$.w�t���"����S���4�^���~��-��&QfLƄH Rw��|*)�J�N#(�F��l���&&!D�VTA�0I�F�t�?`,�ິg%�Uz@E���Z+u��i�~�6�>k�?	GQ����g{E?t�<+�������`�p�<��E|�3F��ʒ�u���tF����[�T��`O�-{�@��)i!�j'`r`�3Q��*�6���rw�Ph/\� �WB�9��:j�l�h䔼$fݬ���6K�\��w�p��ďݥP�����wԁ���Z��0�0�Z2�~#W�y�ԑU�Il�3%�xd���Hd�����艑��Lx�@vҖG�+�뱰�䃗OhY�v����.N2����-Hؽ�>�5��;ǽO�rm�w=O��+�W�=k�J�c���:���[g��&$* *Ŝ��h��r�w�M�**�c<�Qu_h��.�ߓw�S���M��.[���s!�O Z]S�>�\<W�X�R�@%�fsSW�x3�'�O�W��E��Em4����w���#96(�t�6Ь#���G̏Sx��/LDdГ򗸒����sVZ�/�/z�M�x3�/�3�QGb�"�5�K�=�)�����L`�JĊ'�D#��Gg�6�u�LIj����݈2QLn	��-CU5 �(�S�T��?�L���R�t�_��l�Q�^1e/^��L:Ik+����;�c.�02��d�/��� a��^F� �����5��A_�+��'�ɐt_9�^����/)����.�/5��ۯ���ZO��8[l%t�ٰ�O�`nt��4�y�1���)">��F�`�:v4}�iٍKk�#�C�Ma��`?ft&�gdq ΄��������~N�Y� X1P*���nE��o�8mz��1����}w��/�?0C/��*?U��8�c)����~0�`�!��"`(E��՛Mb:�Ջ��3�8ztƤ{졯� �
��E�֝�]�Q�~�%�h���P�S�S�5��s�z�p0� e߸kIe޾:�QR�gpR�.t�<i�Ù}��xe�q��F@��R���!U��<S�' �>g���.���.$�������'^Ic�+�������������g�\��n�в�?杯�P�g�|���<����Ee�{���S^H�t�J����wQa:Y*�0j�ٵ���T?�8JM�Y���P�\2ņ)�B-S���y����JQ�L�o�H�4nd���(�������-�}�4xpΓf�����N����a�[�m��Yg�7i�#ʦ� v�P�@�8��f?�"3�����WB�c�����܌;��Ǩu�4��Zjq<c�՛L9*��m���� �2do��f�|�HY��ܯOf���!׭ߚ�G`��+� �[x|v*�}�>�Wyʈ�2H���'@y�u�%QA�A�*���W�]�b�̮@���[�{Ӟ���A�υ����I�'�XGJ�����nYL�BL��DU�����.}t�=jd��Q��*Aц���ޢ����Ju��aRq$D��NX���8V
$ݺ��ҧ��;��~����l�t��B�Y��]͵�Y&O�|�B�d�m!��Ǻ����/�k�2��"�k��K�,0���w�e�ѷ"� 5qX���o�b�2�E!I�����7SW��L<0h�q��;M1���!䗄EX��o�Gd󁸔��7X��gV�3�5��魅^��[�~h����̨PO3�����>"3bغƠ�� ^'"Po�ϐ+��TVݠ����'B��>� ��y�<���ya��Ю�K`J3wD��ѧ���AvEƅjE��TE�r$�D�Mr��ؼ"�Z����FS;VbԄ�j�yfo�<*GU��Ʀ���.�CZ�U��������c_b C!�L��$X��w���<�n'<�&�x���ET��_��nw���,����v������JV�Y-��P��{���ħ�F��̩�����/.�cI���M�e@�nE��Çb���
>8b�6�.W�GW�ٿ�p��i�����I�	�n-��BB>�lʴ[4M�f�T�����Q�1��ˈU9:^=�^u�����p�]��$Ur`����=�I:���L�.=��!��49�ʧ<��^�v�M���u�����c�(�v�6?s~���r�y��z�-�ԬBa1jy�ˡyU��������Վn/�J���.Ew�aЕ���طWP�~�� w���}���\W�4��s���$���1D͠N��S��*�36��F*&��e��M:F������o|#�CQ���y-H#]R��P:���0����Ԗ(�Lȉ�!��\������t�N��y��E��rtD�!��\�a���J��u���&S��u�#l�!l
#
m���]|3�I Ұ�76p��YL���KVʀU��u8� Д�d�����m���>�Y�ɂ�Q��PɅ��UBV�����9�z��kY�m*�[$�ϼ+0�m�����W@�	Pq���ަ����06$�n�%�B�!㿕';Fo�'����uz��
v��Etl��<�
��L�JVI����@�BF�/�u�`*i����c���m)ٴ"�%9�ãQ���!.�v�j�*�-���y��,X��24-��H����O�W�I����.����uZo���O+�B3qr�h�5��(�nd�ל��F�����6!$�"<�)�F�����>o��(_�,�@Ū�� ��r�0^;�M$ѥ�m��nKY�"gW.-��l��A���=�^Z�>�Z�F1s+E����}��G�"l���"�)���O��!a��E�����/4;b�����is�C*�%Q����X�
��V/�u��C�4�\��\>��B��C�ڔTbqiPm	�dd4t��ZC<!��fX��2#�2�����刲�o,D������H������ynP��f�:���2�a$�ް���H!}ؙ��`oO��j)
����Xۓ7У�2�!�#�o�=M3��-�� ��0��I�? �i;�{�~��D������Y�j.ڄ�=ȷ]�J��ƍw��[�;�{��`I���w��=#����w|����0�Ծ����<���0F�4�Os��\v�n�Ky��-
�Kv�Z��#/�� F�<�_���&�%GO>�a?kI�o�������`z�S1�x?���l�F��J^�/�=9�e���D�P�g=Qx�;�{Z���q��~��S�r�S�~tt��[����1*#-d�7�����&�B�_�'fܰ�nr�Ex�O�ہ�z����1>��͹��˕�?H�`��������<�ٟ'z|^���dW��FohC[߲/*][_��d׃IR�F�v���� 8.�b�1%F@��W@�on �H�.]+:��Q��FĪ�j�w%�����i���E�lJr�	�~�Q��<}ǮVdՀ���~��Ä��U-l��bn����q�`sP�d���	-�I��PO�B�QWt�����Z�������u �.eAG6����X���������S�wx�=>��)���x6���b�HW�r6�̡亊��ɶQ!`I��D݃���=�e�|��#}d�����M��R�䕼��q⚱46�-P�ѡjA	�fD���8c���,ǵ2^F}�̿CMr��탣tG�s�&��H�yi�M�Z�T�Cf�΍��Q�w �9B����ﺘU^@ )�Ҩ�#Һ?�L���ڏu��5nY𤩿[�ŵ�ݥ����`F'��/>^q�y�?���q�n�`���;��+<;���q)�(���z>5E]����9뺱s�L�H���E��#\�qꍰO��
�Tk��{��D>�: {{E�eG
Z,�����һ�����?�s,�h�U�վ�Fׁ�%���=�����n~+P���i��Z�lׇ�M�*9ʹԩ��.��%�YmW�S�T��ǝ�IP�,�6�3���O�1�c���?0�f=L�X����D*�R�uj�u���\�E��t�ϐ��W�<m&jޚǒ_���"�W�7;��D�h��{��������
I��<3�bn(C�!` ��_ᜀ9X�� _V�J���p-'�G�ks���Y��a��N�����a�`3�T��}s1X�e� �0(�9,��K����ڴ+�D4a{����3�|��)n�q'�aPس��-5�p�u�-%r�O7����]� �.��5j���{4�y�K�����^����v]���O�:���ۨy�5I�W���(�t�g%V\����X�FN=-9���ޅ�\ӄ���J裸q�m[7��-)��B3b�?�`�J�Cmd���x�.2!��&�Fd�n̅Ku=?�l�&�c��Έ��>%b]�%��<���X
T��;���N���z�?�/�~�-�Yw���r���Ed� F1.��|�ͱ�&�p���8�a��S7���U�=Qp�q�#J��a�w����:sI$*�����Y6]���Id맟�k����{s
���h9��։�i@i9S)D�̬��gDBr��c�[�a��F]2���On�G��W�=�6�Be�����r���䒮���(?y�h����L������+8�|�����'���+��o�I@��{"����߁�6�05�k-1s�J'd�U�@�J�ʹ��\իE����	�t����S/�gU򱊝'w-�Gm����v�[�|VW3���4�]��q��Y1 Hd����^���l��KE�a�ة�)���t���(�%n�5����8��ƫ+ߠyٿ?k1�2I����p?����t�F���3��_d���t2ٍz��M��d[��ƕ	�Wc)�짝�u�r�*�S�%�;m�S����[>�ruB�l�W�\��\4Wާ�Ʒ�*�'5Q+�, ��`ÃԌi���	���O"�����gh��7�B{��;��"��� ���_`c��߳U���r<��I��K�.>��Zt��4��i�֨`)qHƎ��*-�-V梃�ah㩞�d�����Ph.w�(���<T�fRq�S�O�l����(砒�hC2 �����	� \[ڪx�g4D8g�� :�L�'��lĂ�qF�`}�W��,.Vk6��x�W�'��1�2J���C=3{�����c�x�)1�46D���*h,άk-�Ԃ�0[V�H�,���p� ��W��=���'.��uA0��rf)"7����G�D��1|n��Ð]̊$�yH?�ex�Ju8��|F���H��G��&�� 4Igi�#4���PV�6��U��P>3)�Zӑ-L\k}��7��V~0�0	�y�TT	N��6�7�c��v��WI/	�L�OH-i~Xu����!�ŧ���_4�\S�{�~���w�g2
���W���J�L���񌠸��-�%��;�l�
��X{�j���J��Yp�߲�5cz�|�P���ym1�� '��+����܂��	L���ѧ�MW��Eȯ��h�`���uN��J
4��U�Vx+ڻr����o>*W��Le�KT�q�������+Ȼl�?����9?�%x��t�@�3D$�b�Q��hB�����6%cV���	�t�!m��� ����r�����m���/�pk���!�25�l�)sc�(kcD��w6w|"�m9�=��h4��Cx��X�NY.K��TD��)����rˤ��u.��� ?Ŕ�>%-�gthm�l��ǨBB��^.��^+��	�!��g�����"3we�����+��4c�����|��`w&�tD���FsT���c#}��1��\w�6Q��e�
�P���l�m���!OPhc��װ�Ǚ�G�= ��20n1��k2\E߷��$N!)�B���잖%
;����@��j�����r�֛et)�r�tː��H�ѯ������{%�ᑑ.J���c+�+��nn��D�X�-��ݠ�!,vC��\틉�K;i�Y���D+*�0��dz�J��D�@k���G���%+c�<L�HfY^����q@���f�9'huܣ3m�I��S99�p��^P�v�����-��6���%����5����{�ڕ���h�����W�8n��nu!��=��!���=_��8�D�]��u[�r�� ���:w��Dg�w�8]���/��}Z���|ɂ�х˼�F��VFM�·0�X�3N�{�!����j%� k\���|��A�@L�Y��Ԃb���KM��;�!q��kn6#����I`8�Z�S���4#f	��	�]a)��YfF� *���7����`��?ٞ.�\|M/�J�w�������,����~х�u,j�NK�����	��Ͽ�Ȅ=�f���u.��'�.a���C*�2y=Ԍ�yf��v0��zɭ3"C�T�d8�Fe�6(y��4I�����^6d�+��cv�Y�.O�h��wt�\.$��8 �_�Xrc5���^^�;O�`��Y�y�A"�}��8�̌�X-&VA��O�sX��v�:�z��|9���3��O_H���y�V�ɿ4⎱B��èչt5�m���Ә��?r�55��ʫ�Ѧϓ�x����6��`�FM��6���xL����pO3��p�~M
e�����\�:uT=�9[�v��e�+��1�;V�O���®͇	����x%Ϻ� =��F��`��*z*��@��hf(��m�bm�����(�l|��ú.ʑ�G�����O/���vv���"�����)8Zl|#,�/��Wܵ�"�{ޝ&LW��#a�9 ڐ"ɬ����ŵ�j��YW���l�^-�y]�a@6ĥ�6�t
'���vu8�h��DG���^!?9��N��YD��n�;�6�pi,EV�MٝW�b��c��O����JR�.]��V�1F�YA֙�p3�H�^�X:�9D�7D�X���\�%�O1��h�$�P��ޚ�6�Ns��6����Wq��渻�]��:����MI\��@~���]������:]���Q-�y�Mi��4o����!�{t�����t����@`��ߺc�c��s:��	�֒��e���=/�3�3b�
M��ӈ�57)|��q�
�
�]�e0�R�r-�`�]ˠ)I��JE�g���{){��)��P��ʘ����6�TI�������� p-*=M��Gl�]q��S�Ҵ����I��"�	��w_���t��L�:����@�����r�!"����$A���D7O�628{1yu�" �г��H�gg�mgJ�'���}�a}��2����J�:I�G?�C]�bB��1<��f0�9��]�S�S����5E|��b��/T ��bߥ��~W����ص}�n ��=�0�W�<c�n���s�9-cBDf㒁�+ܓ�J���1�*���
W~�6˿��eԗ-VRY���)�ơ��~�ADW,���f����
�̦>o�
MPX��^��liW-+]?󧸝`��f#�;T@��5�I:b4�G�еk���'�R`GQ�MueU�mќ��ې��`W�Te.�)�%�������K$��0�\��3�ч�޳>�z�G��?j�^)V�TJ&ן����
�r��`.��e&@�|l�)�v'��@j���=�ĵ&c��+}(��y�SdZ��9������! v�%�:3�.��7u���,nE�z����͞g���ג��L��9���~<ћ�pB� _��=���9)�������~}ޗ<ܱ�!�<o~ªnW��t9����F�G(e��͍|M�jl���zy{"�+_7�kАF����-�@n���fT.��K��o=�I�'����x�����n+�xT��7"4�M����00#U<��c�2��%&D��lx&��`%5f9#��&h�5��`6���㩜�� ��
M�op���:�j��0Ǜ���;@L���pi@86����q=�n�	"����g̓��V����o����B���j������������!�-��Jƃ�^�:-�x��O� ���T��QZ�/Y�����ձ���	Q?�BP�p�����[������9].��6�@�O!I��f����-#4�a���*p�:jMw�v��Ļ³i=�z�9l8����L�����4��Ob��k��z�a��`�\���@Z� ���n�,��^zܧ�Wk$ED��r[H2�Fitj����]�%J���u��ө	#bxdf�m7�~�J����$	���T$���B��ܤ��t��6fs����f-5[��&��7����HU���mݚ��<�+L+�� Խ�t�֦ϛ�EmGǺW;�1�d�a��/έ�޶T��6�X� =��m�
q4�t$����Rמ�B��ĞUi��Y���ڹ����$?�zĠ���6�_��*ۨ;c��m/��GP��)�U��)KzҶa�k�����n���E���N���Z�4բ���e>S�YŜ�s���3c�Ł����KU2�Ui�8�v��v�l�吝/?��~{��KϮ����i�Lh����yN��s�#b�H��ꕖ(~	0oP�gl��|�p&��E��<XĿ�ɠ�9>%}�R��O�.�\K�0s�r^�{>U�)!�T�?����1m<�v�h;q���!���r���S`��$���Í�8J���Y���I ����e�?)��[8�;h|�Xsb�zyc��/�����Oy�̸|g�����Ҹ��3e� :4KV�]UyY/�No�sQ�^Yy�U�%֙�%E}�L��PI�;�H�|Y@2��3&:�Z�z?�2�,JF��مK�E�# %��~ۜ�4�F;-~�B!�nHޒ���HkU��>{�X��6�/n��E˕<�yͤ��ZvV�A�O�H�7�&����(m��(��,'k���t�L�y4�d#o�P��x>`���.u%?�<[�����
"�)O]���Ž����mZ�C�-�&��i���5I��RA�	<�o���ӛ�Q>�<n<?�3���9���R1B2�4�3��mf�!���`�'�g�}���s���p̪@�	��S���rH~�B��2K�Z�]շX��ZdY`>�$	�~�zm�]�+���-�	����6�W"�lԃ=��j`ν��z#�������(�u���&����$RD�-Ⱥ���ۗ����^(@�]}Gت��r�kj�������jI���H� y(�n�h*�3j�Ίю�AB�(�wz�p��jf��$q�"	�W巼o�栞�)Z�7�N�a�ǝ�Y���=X���e���bW�����I^l�3��ߣƭ�����߀_Y1��2��.��Z<[�'ܴ�U%v�� �:aYKW�xu�����u��Ŭ$a��V�T�k~��=u�l��&��/�3�����kPn«6���˻�p�@��Ņ+���V�=ȋً&d�����:/k��z���~Tqh9�R�0�ԫM� �f0v5B�˷���v{���LzX�q��Vu�bZ�����¾��ǝ�/Üyl\���+�.�<����G��"��y�O}�ZQ�B�d-��@$,T�w��s��
�j͢pz�Q�MDY�_�*�3�\V�)ad�5�]a����"ts�3��܌��s�_���i�	��c�>�t::�`e+��L^p$�Ǣ1����w4�(�A�O21G��	g��V/��L�]!�ȃ-g�G���������C�
�{�j;�O]L/�-��b�[^�j���K��Ʋn f@�$;�o��y�������܇y���V��m8����M?�!@�d�[����ڗ>>Mto^<��=6��*���Z�z]�1	�j*�`R?ـz�B�A��r�s_��_�]��j)�[�G��T��W��-!}b�.����,M�����~G�K�$�Ts������-a��tk���A/��]*7�n���y������.ô�۾o�p�0�I?��Ʈ-�����n��.g�i�q���&�z�tվ{�-���{=k��W~�3Q�	op=���`
[��ƃ5X�ւn���?Fs��Oփ��y��7p6��Pg�?w�0���G��iϻǥh���}��Z�V� g�.Xu:K��������Y�����P�A�ga��{�د:���2xE��l���3-�� U�L[�E�v)A�,5�c�r���S���K�"�!k�}�0(P�lM^��M|�uf�lip�ݼ�}��MQ8O��Ԣ�S��B�w�~}ou��H�Ioc�u5�z�������m�ɟǊ����o+��ؤ=��!-|4w1����U�`�qBx�=��t�5ϙ���J���^Cdf�����O��h@@�7�`��9=>r�!4���;&����|V%�m�&�KP��8dm���G������2���j&��,�D�5%M�B�rO�F�E��k��J�P���qq�t�9�BQXٻ���I�wd(�0�u�<�����u���V4�E��	#�хs�Y	N�n��4�IVY��3�7�d�����%M����c�"�8P�2��T6��Ɛ�\]o�_!]0M�B��V�>�� qr�_�HW}�US���o��y�[lp���@!p��[��q��t񋜑��g�j?{��<�?ؑ�x	�e��&��ϗ��n�]<�R��(:��Vrp�!7�X�^��ʗ{Y�e���X��=>tY��cL�N3�L����ЏS{l���3W,�Wj��ځ���ؕpDU���,	Q�L]{+��Z�cL	�0�s�k��:���$���Rk^b�%x��Լ7��������*�g���S��i���eVMz�h	�">���		H���N�&���f�nm�@:LF��Q�~q��gL�F��3Y(����Y\�q�U%�rnp�� �(=�T�T�H�]��C젶�y��`�&y�����0i�Hʾ���h����᜴0�e��2ꂊjQ 9n*K���EhD�spE9[%r�	V�8��%+�Y�i=�{i�����{-*v�ߠ���Z����
)��#�54!%�.����l�����ǟ�S8��K񽄪*^;�W#�P�S�;+�?�iQ�l�F��%6�ŃߔO߫T3��,2>�l��%��ߥ[�iK�K&�k�1$H�$#��GA���O�'}����~�K������7N������rX������՗k��i#vR ��8� }����{���%eo���_��HV��°��-gY�"Ze�$ݵ����s�/H�H��%C���7�,mc����CK���PP[i[�9)�s�I����v�wA�h����[�AE���"
d�f�.k�&>�a6�O������	*�_��`+��R]�KƏ��\�ઘ���u�j��r)Yh�d���<>���;}@.
��t��岐���L��4m(?��W��h�N����D��>����?�&?�sمf4ŕ~�C�_�3;w&/݈�q���ζ°�}�f�\��Ͷ�]u]�n���FZ�5��������d�����{�KX��~[����T;Zߧ�{o/����((�aƚJ����@��Ӻ�Rh��&Nz[��X��L����T�*��#t��}\`�3[@	�����|AQ����VW!��F�~DH�2XN�'X�Ԇ'�������w�&��zff3�*Q�P}�6�lk��E����1|"|����Xa}czļjt���S���F�>l�>e3��^��ch�0W79��n�.�A���S�+����|��a��Ɲ� 7�L
C�d-o�\���w�PZM��Rj����76�Y�ww]L)_/
����숒y��9��om]:�!F��N��ә&�R!&����N�Q�b {V�2�?�@�IHN8��0{��qU8F��#n���\���"H+��᫇3xhd>�k�B|֟^��ɉ����f�`�yHBU
�m��V%[���Bv=;�t�G�C}�W	����	3�'�@5�6Rr�78��}I�Y>?� 	�+�)I�*�O�
4���B���@𣐷:&��<Ka���L%G�?���J�,����E�#4n+���9��t�^���L��@k�Փw���k�	��Y�ϔ������MA��:�k��r*�}���;��W�u�:7��V2�]ē���8����U�Et:G��'5+~���0�H�+� J}���@ti�`��iy��%��s*v�������G�պWt	ϙ�ݶ[M�xJ�;��xZ� ����ޣ�M�lj�2��{g%b�2�` �i�vPc]'W�nZ��1V�+��a�,0<�bD�D�H�{��M�u���F���puLN�8��;�^B�C��!��Ǖ��Nh��#Mc��jE���JU�����o��,�ʆ��_����~��Z4*�Y�<<c����)o"��8��B�� ����{59���Ǘ�t�����T�g䊭���	��.�QOe������PhK�FJ���i8�@�E�##��Z�_��02_j2s
4ΟO�����_���v�_O>��⒀�O�wy{Rn�z9f�@�t9c��W+��2]�K���m��/U�w@9ވ�;�:�3�]�mg���Ϳ�����8a�C�R9�!��j��������gzӷ���i�l�S	���Wj��Q(T�2W��}9��\�E��pЮ0|8OE���3������u�65�M8U�
Z�?{$tXh}�v�{[�� y�3��&���m��,�nL�������f"�eKqQ�B>��Q������6Y�4��,�\K����#�o�����}�xbFQ5���ј��R*8��O'�"�����e`
��M�M�ԕ�=�	�_���5���;���#/;�aN��4����sL�򚰤e��Fz���n����^�#/g���`�W��({�3�H�Yx ���5��L�~X��D�=�+����R�%G�X_�~&�'U�مX�(�q�d�sp����i�x3k%~&�AD���,z��Q�
�m�I�a��ZŒ�TP��]���4�C�o�� 7g�*����,֟�S�:�����n��a%)�6?I���>;�GY��u؛��g+� :QW28�����-����c�6�Ӟ����>g�T��+��my��!��M�y�7��5s5A0���9��Z�ś��
%��"F�17Qd��F��˓�J��8O�iaI���%nh�cݪ����<�'�J��u��-�p$� 
�5��:\��o��s�('\쏒�@d�־݃�ֵ�YI��5섔�kEJ'��KU`4���P�b0�� �1�u�J�E�c�Ïh���NN�)Ӳ> �<�+ ���[�Z(���,�x�-Wd\'&v Ű�����F ��H��;?��Ė%:�\I=��/�=�B���6��[[VC{�b� J��h��mv��="�/$�MAVUfl�e�U��0�N�H �3�"Ss��I�}Yr�۶d�4�7�����\���W�tb�G&rk�|fL��DL��Lq:)e�m�mm���|�-��BQ�4{N�ϩ�Qq	��\.�^:#���5o��4ы��Ʌ�C�S�̄8R�F$XJ�ǵX��2�֯A��YIc�K+�}�rf�V��ؘ�SBm=�$�������P����`��փJ�^�~B�"FTw�aub3��U��9W:.�5�@���*G6�^�����;~�R/��Sa�����>��J��iI -���ҳ. s�k����E2�����Y�2�W��-.�ACS����C�QJY��ȨhZ6~�V�M��5���ҕE�9��v�؞�Fq�f~�����]�ߵ�2GMf4��J��CX��z��W��*�.�jN\����jq�M�;��{��몕P��K�C?�@GJ��x|v2�f��h�t���m%/��P5.���N�Է�nG��Ǜ��ޭ���A�����w�u^b�}��tp*[rT���C�Q)C�M�u5.sh�}x!�ϳ�S�c���'��U����آ�r�t*�M%x�裢��s.��X�n���)�=��w���P�əC#x�Bg�+�?����Q�U�l}�L�<���͓?�� �%�kԋ���t�ƟuR�љ����G|���[�O+��0�a�d�*�jr�(�M�.��2V�� �~���X�?~7x�fɾi:����|IO'�J�o�{��z":찙d���f�/�a��7�& ��A��>��y�n�'Y\�e ��ؖۘd@B'	*/Ou|���=�O��_�@�ZU;o��r/jċ�����v+}Kȧ�c)��`��o ��_2�����ٰ"�j�w��Y�A,�\?�|�q�sՄ��d�\6.s�w3Ss.z��{M���L�ߤ�d�yZ1���W7m�.���|�ڜ�=���+�G~�Y�3��|�+����7�z��e�҂��c.��=����L`��_B�w�'�W��m*M6��x�Y�>ɊeO����,���Ɩ�dt�̛�'i1Y����3�O$O�(s���?�����_^~�7Q�h.U�4��>�E�|�P���:=m��n��I��#��������:��������X^ 1N�u�)`q(Ur*2D�P��p��p8��}�*7}6��|sV.�����S$�=�sn��	�b��=�ޓ�%��YW�J>�v�&Kd�BmL�Y%mkM��!,|vKȄ�� '�3��ў*�@���)���^�񖿡�<�Jl\��%��<Ts �ؙ��h�[�(Y�� -2�NR��S"i���@�MI�U�̕2�F{�,�e�&��
R���Q��� �W?��M��M��TV�w֌����9᭪���	�e��?�u����Rt�Ļ벤�b��1L�q�,�������rp��Kh}��契oʯ��1�kH��s� S^���׿��B�^2_I�����O���v7�5�J߁SH��E���Q�l����B!Q����΄0����כ~����<'���Ǡ7��1��R�O��x�ގ ����. X�N�О�%i����uF��D�!����P�ˬ!ܾ��z�k�^u�K��������J9�)''��o��%9u`���?�Cy@�/���15�:�.:S	4�S�r�7}����P_p� �{�O��}Ty�$c6��(j��Y�R�ʔ�n�*I���P�m�>WsH k-�	���i�D�1��@��AȦ�e$db��	�3l�<��D_���p&�5(�<���"�;��o��=I�*q�Ë��bA�B�~�;�;ݦU�S�#��O7D��DŞ k����**���
3l#�|x�3�P�%/k\�X���|d+�J֜Ҽ����_2��I�m6�~W4��E�j�Z�׿�������|�}j�l0��k'{.��1��B��~�i��kL$\]���4�˅�	�皇y�^
4Į�R$Q,�B�2���2ֱ���3��
�I U$gتQQKU�F�m*K���a��:��,8I�C��e��2�Y؝C<�48��Q-Ձ��۬��S3�(�uꎊR�*Ik�5�?E�Ҟ��[�ǹ Y�]���;lPQ��I Dr�)~O��D�{C��^�@�ە� kd��*��狡v� N�ԕ��n{FleB�<�@��i°�����i3Z̨�m/�oa�R��������1�D��s��t�؅l'~��m��k���|+ �mV���נ�>|���]R��+�I��4�j!g���[�����:��2��b��;�d�-��� �^"��6l���A3��ý�m��&�7���&������w�k;��8��b���t��bx���ʨ0���E��E"y��f�hُ���B[�h&�����1�o픢^�as��`p��(�z��@HK��W-p�[�Za�qv��6w)��^�) �b�� �[�RR��F�N�~3��CUǕ�=��s5t���b�\P"#b[u}kq��x�%��w�i��콚h�z=�� �M���F��a!8"?�lM����$6>��p�0i\�N��[�s~5���A������@��a��h����;�"G��$�R���x����Y �	A����#��L���)�X�����Ek�$���pƸ�X��>�7;U�T��Ox�a5Փ�|q����$��}�(Nu��à��-�X]���{������C)%����4����'���ʄPpW�����8��B��ϡ&z���yZb���L"���J��4���.�S��1o ��s�x��<Q��&yћ�fy<�)����Q�p�����-~篭FxY�A���q�n�������H�3r��Xs%�.����&�CN]O�_c㌏~�C��X#q��!�3<�L�N"�dﲻ�D�!U)>Q��M���$�
�OH0R$�?̘�d"t�I�e���]ι���V�a�%W���_��#��;�>�gԺ���[s������p�bD�t�'B�Q�yi�T+O�C�/�HId��,�����w���^�����A3��s�6<U�8-���P�rva�T�<q$S��h�+�7���L��X�nz�a��p<���F�Dd�,Jl�{i�>�4%y��a����~(3P���2���9��|�"�M���=rG�|�MN=�����V�HLj嗶Q�b̠��u1�x�>�"�W��/#+L�FX&6\�󮁲�Ӭ¸���.����&pݕ�G�3�V����D5"m�9�`K��D�8��\�h��u��w}|�y�,�=}���'
*N�S�����wv�%���U����#�#J�9�L�e��S�ۡ`�$��'��+�6���k��w������+��	��;��
�)�x�2d�Ԗ��fhI&p3;����f�ɆJ�4�_��hS��	�W�������J�������#�׮F�K�B`!{�|�V�Z��c�<��|Kz�E�<)q��&X��Do|���͸Fɏ�R}����5�qS��˴K�R(��tR0���P&�S�-���ڗ��:�֒���u��a�i6���ϻ>^�Fy.��,��]c���^�*� Y����v���9c�-��)���=�(�,���C�b��e��`=ޝ������#��L�Y3����Q�����p�z�;4�������I��|����-v<�>d�w�o`�b� �w�V:L��XF�x�
��Б̩I�K�PpD��D� 
������k0��(��Q�,x.�s#����L�]U�O�F�R�Y�M��7��{����65x�}� n������!�����s��	��o�l�8W~x4�S��Y@iB�gN4�t��BB��7���f�nr�$��A��x�9�/�T��W�R1���`؞i@��?ơ|��_7NDm@�1Yf!��Ϟp�Q�1��Jk/z�^u�?;���`�p�*�/^]	��~E��-�Ɠ~+�# ����9m<�;�h�����X�G턉qȵ�	b%���l�������ض��{�Z(���]S�]ث�ˠ����j�
{W�ILU�*��h�؈JA�R�Ր��Lt��7 !u6������߬&���O7�׳�G�0����.�g1�e���J2�{w����gve�5��.4��"�	�},��-د	���pM�vۡ�hљx�9GLLsj��B���rCy�l-+������W��2|���<s���T:R��
�x��Wd�b��4�fW��WSD�e�J��t
C	9�>�B��Ji��o`�~Z2�bE�IC���R�;<�Y�7��(6I��[;?:�;�^Z�C�S@X�6.���|��V01�ü� N7}V>�����Ȩ�2}I56�Ż@������l`j������ge9�Y�nf4�-3\�h�4�2,Z#.��`,���:�8Ÿ�%YT�@D߲�X{�2����ЏE0�e�:�s?��d�y"2C�3�KQ{��c�tu��E6ت����ƛW�{��M�t�W��	����x��h�m��+��ޖɕ q�_�( �hS�	���A\���6��\]�
�� �ԥ�2�Ѕ<�������ѿpߊ٪��P��RxQ�R��n@��pv����
��c7��<C:6�׏�Z�D�s�ӸX��"}b�8�=W�}��i���t��V�7�W�2	J��Le	xN�����P���&rqQ�����UK�s2\���x��:��0�L��5�&� ��r)�(�l2��!!��/����(���CKH��߽j�cc�3bG�n�����i���_�Fu��J6���B�zXwp�����Ms���(�3L�XL�������-Xo��z��x"����'��T<X�;�rT0�ύs������crۆݍ���xa�f8���1��z"s	,�D?X��~-�\\%y�_qÕq��}98jw�����D�����w|>J*RZ,�y�r�M@?����zz�U������#Ů�б���=��#�!����H���eyI��C��ʅ4��{���aL�E).�W�t��չ�
=�����=r�t�%@��42 #���\�x�oCV8����Ϟ���g��7_ĥ�k�n�~r�.*�Ms��y@��������w��md��s����b�+pF�E���������7J��M�v?����l���^�L��F�*��`xR~MTF:e�b���\��i�~<�����=t`�k���̸|�s��7��d���5�bQ�eI#q2�߲ի���_�1�/J�[5Y-�)�2�v}����\ ��i��N��c7������^
�N��|����;sE�Z
w�
Y��nޡ�m;�"S��[V��zEv�ӆ���r�O�˓Ht����Mv�/��0ցx�����@�[v3�́��;�N	� 6W�@������7��΁�SI�g!�sC?�O9�Xg�1&�3s��J�,n�'<V�^k���ɬk�b��R�sa}�{�jf��nhZ�y�~�2�j*�J3t�� �:�-.�Ĵȩ4��w�1'�&h!���G�5�ɾ&ș�l�+=�&>rE:�c6�)��W�d����ׁ�-zQ��>�d0n�Hh��$��	!��-�B��:�:m�L���ˤ����SO�� W$�����_ƣ��Ǣj.��`�f��@O>n�źY?ʰY��$Q��%q=2���+�I��y*g��jAdj����އOr0&�#0pA�D���܇m��VA@��p'�Us��y��ku��~�F�d�,>f��ի<&<�,��6ڰ�RR�x�OB�s�]��`�t��z��q�d����i�<e@�y�9D1��.�|�5x�Dx�"�8/�{x�/�ZFNoE��V�M�5���A�����)����M�0�\d�׻Ty��`���b\�mI�yN�ARF�|�]��M8v���1��|g&����]�n�U�?|��3�zp%m4g��R�4
�'S�E��Y�~P%� �=�N����ѹ���u&B�Ò���^_3�0��%C^�
�l����/�6q���J�O��ן�{z�6+KW"D2�6�WlW��1-�&c��^��i�LU��z�9�Jt|O�.�#�Z�M���_��@ �Hctn�4��Eh|O� =�ȅ��%���r�nh��bVl6����f.�?��I6C�����DY#`2�8=��z��e������`WV���O�d,ٔ��Ԝ������3��r���cO��1��+#�Xt�0��8�Z5�>�Q�)K��I��k�$��qAVo̇�vj�1��#\i�*��p�r\�c�Z&�9����7�\C�����^�{�6�)�<8���
6��h�[ż�εY���l�}�.O#��M�6�"�m�e�,:�S�L�[��Ծ�������v��Ǣ�g%N꩔*t�c��8h����t7���ϻg�Q���3�����j�w�,��cJ�.�ݢ��_#�s�t���PF���?l���<�1Fy�Ɂ<�����.r���nϳ�f&,���Ү
��.���r4:�W&U�"m�h�g��ɁP���} /ļ��Y��F-B,��K?�oh-�*�H	S���T:��z^(:&
�s��� �Y��5���ѭ�M����x�Kx~:6
g���M�p���_�V��%{?DU��ဩ.�c�����vnh�ē�`1:���ҳ[&���LcP���fm�K�x�����Z�:�4��B/qw�T��+���mK���V��q4�t�S瞗xH�뮒��L���QD��͓KbC�8�6Z�0���=0/0 �i���NnD�A34i�Ew��N��8�K�`��"&Xq\���?ڿښ�� 7�a`dٵ�x�7\(��Ce���WrJ��,����'a �D�)̐��#l�
M�7{���S��|u��)o]
jZ���Z�W�����@$e$��t���+�P!ŝ��ճ�J���M&��Zㅎ�3�@�/1�h�����K�0k�ec�D��ƨh?��8�5��#Kb�1nI
II�S�:s��՜�Q��� �ϑ��""*��KG��Ao��~J��Z�Y����0��:1������N`\���՛*���"?�`��_���e|��8Ḷ�x�#�Y��=��~x��Y[�+KO�dB��Mx�xa�o���b����9�0�ۥw8���l����>~q��I����_��1��`k�)��a
��Ĺ�0]E�[���1�;��1�"F­!ցc��ـI��=�|$��	<ݛGh�S����~Fct�`��T��p ^"n�3'��	��/7A�j�x$_��p%Yh�H�^��%�I��4�@��|��S�P�Ro��P)�Ч���R�"s�\���'RiN��C���!\�����,��䫲h"񏬡
����YUt_�� |e=ÕԌd��8��%OD������<�My/]� �h�xw<�قDm#���ZD����	L�Q"�J�K �My7a��+�
��Oۋ�����VI���kK����S�t��g�Z�e���Q�
2G.���<ᗼ̻�����^'ដ8:�JB��k9f�ɸ��f�������d9���J��ܺ�7?3ޏE�$%�NY'�d~�S<�+���rR�pl�1�ƪ�e���8}���"v�&������2�������]�q��Q�8I�,��B�e�q�Պ=�}��EN�>d��*�d��8C��Y��J�#�B ˃+��0\��J߲L	�^.��^��n�b�:>ڇv�߫���2��	8�V��i�n����s�x51�-���i�*���*Ye�2��ɓ��M�6��&XBj�o�I��2�>F+uj��Z�Ӧ�ˣ�����U�B�f� �A�o"�?w�
��<�!ގ�̤���Ӧ�-i?����x���4p�?3ů�D��r������(�~,�w�1dO��7������=��(&��C��G�H����aB��cy;ƞ6R~�6�(�a�j#s��t	,t�@��ǌC/Z`l�J�E�,�7ִ�4�-tF���i�t����Ö_�� ��K��ӓ�z�S�*G4�F=o/�tR�P�Bb�텲��9K�j��xO�(�����3�p���UL��uv}�#6�I[
-�z5��B}��7�˵���脰JQ�^7Z.�.���~g��� U%�����r=�����9IlG��dbI��݂���ߦV��|; ���^]Wc��"�4i�e�Q�����er������ 
5͐r�.$n߃o��-^IN��"X*����
�y�{���,նn8��������9�	�ټ�5�k�g�i�Z�}��)���ĻX��	c���<0Y�*��z�8ε�Q���Ȉ���� ���Dd|ԋ�di.B<��Յ��	����ۙ�;�+�ǣ'�2�V�ړ����[� 5^Y���3{4�Ó�;�#|�֤�e&1{�,O����:~��b%=���z ��ϐ|�N1%��6,�8�,�ц��ƻ�j��|x!h6�S#S!=p�K�Ү!�w��&�ݵ�T�����|��n*K���(S\��	+Lck�U[����2Ւ��@�M�Yτ���5*de�_bk�2_&��lW�C�g}`���$�7!��9�� ���
������d+����1�0�!_�v�3I��S0�Q"�*"�v�d|HԻ;'�GLG�5�S�r���}�]�d�b��}����������	_`.�u�s]S��rz�|E���Ə�� *�!�/sV�o3�\�77��E.95���9`Q�<F�s�o�x �в���ٛ�E��2��v�����q��Eԧ�߱��E�����d�f�k��~ͮ���J��WA�n��.�s#�1	xj��%/~e��!���:�� �Y]�*˃l�����Z�Qy�G�Ј��"U����zX"�f��P���tP[�����9�r����a�续��
��CzyH�����pRx��9���Jh��z�n��|I���a$kE��-4 K ��ݏ�~���%fy�.
S$�}���&&��*sC8#���Y�)����P�ҰD>�4�C5���`��:��})���([ ZD�,
�L��6'���T�!���W{$T��!\M�Vd�S�h��ocs�4ĽN`�����0����9	���T
�zV�.�-M9�y�}��!�
/��љ�B��.J�f]�S���ם�e��d���ea��ڄw�N�o��=S>!łE�tϬ�T���(B�֏���.�rühU��,2it���!~�?�jl@�A�T$�`^� �:�?��?8/�l}<��[Gd����;j%L]�n|Fְ��R����Q�c;���R�8�b>��n`�T�}�!Lsx
��h��뢴��Q,�R��ʟ4�E� \���k����X���X�$�q��a��G�W@ю
{rW!?�ϣ�,疏�g����r7��ןכ��X8���%C�>8x(F~�N�]�1�x�[���0�ۋ�
^ד��=)Pc�	,J���� r���Wf�����Ҕ/v�����,0���,r��_d=m�~ �wj(;�
��A��q9�@�ѥ��s��V?�p9���^�|<ΪK�$�1�rlʐL�2�t�[���GGFv���7HG_ِF�#������t߆	ѧ�������%��N,��-�RP�G*�8JB~���@t�Ѓ��C&�����V�5d�쫎	������H�*w��9��Ou?+&t�N"��� ��)��C#�."6Xm����:����35���W2�����
(���jy�P/U�4�����iM��'�5v��Ī�g���a��0�f:h}pnM~$'o���?�6~�=J�I�b��XE�^�@m�0�<o�trz��hk�ne�GQ<A�+&Jm=����%��%��%h�z˯{r�%=�� M���r©���������{�e��	���<o�#�K��d�u&�N<ImdzM��7u�a�j|]_�����k��SO�V�{��F��11�N����y��v�寪͆�(C����c�*LȴV��R���&�@��#�AP�%&�~o����%��j/#������da`���O����č���:�Y|�ř(d�A  �Y�djo|��y����O�60ӡ~>�vW$�=9}�	$/�Q���hrM3�O\Q�V��8=���